
module g07Arbitrator ( \c1.sysClk , \c1.Breset , \m0.need , \m0.ack , 
        \m0.addrM64 , \m0.DoutM , \m0.MinData , \m0.Tdone_mstr , \s0.addr , 
        \s0.SbusIn , \s0.dbus_out , \s0.en , \s0.Tdone , \m1.need , \m1.ack , 
        \m1.addrM64 , \m1.DoutM , \m1.MinData , \m1.Tdone_mstr , \s1.addr , 
        \s1.SbusIn , \s1.dbus_out , \s1.en , \s1.Tdone , \m2.need , \m2.ack , 
        \m2.addrM64 , \m2.DoutM , \m2.MinData , \m2.Tdone_mstr , \s2.addr , 
        \s2.SbusIn , \s2.dbus_out , \s2.en , \s2.Tdone , \m3.need , \m3.ack , 
        \m3.addrM64 , \m3.DoutM , \m3.MinData , \m3.Tdone_mstr , \s3.addr , 
        \s3.SbusIn , \s3.dbus_out , \s3.en , \s3.Tdone , \m4.need , \m4.ack , 
        \m4.addrM64 , \m4.DoutM , \m4.MinData , \m4.Tdone_mstr , \s4.addr , 
        \s4.SbusIn , \s4.dbus_out , \s4.en , \s4.Tdone , \m5.need , \m5.ack , 
        \m5.addrM64 , \m5.DoutM , \m5.MinData , \m5.Tdone_mstr , \s5.addr , 
        \s5.SbusIn , \s5.dbus_out , \s5.en , \s5.Tdone , \m6.need , \m6.ack , 
        \m6.addrM64 , \m6.DoutM , \m6.MinData , \m6.Tdone_mstr , \s6.addr , 
        \s6.SbusIn , \s6.dbus_out , \s6.en , \s6.Tdone , \s7.addr , 
        \s7.SbusIn , \s7.dbus_out , \s7.en , \s7.Tdone , \s8.addr , 
        \s8.SbusIn , \s8.dbus_out , \s8.en , \s8.Tdone , \s9.addr , 
        \s9.SbusIn , \s9.dbus_out , \s9.en , \s9.Tdone , \s10.addr , 
        \s10.SbusIn , \s10.dbus_out , \s10.en , \s10.Tdone , \s11.addr , 
        \s11.SbusIn , \s11.dbus_out , \s11.en , \s11.Tdone , \s12.addr , 
        \s12.SbusIn , \s12.dbus_out , \s12.en , \s12.Tdone , \s13.addr , 
        \s13.SbusIn , \s13.dbus_out , \s13.en , \s13.Tdone , \s14.addr , 
        \s14.SbusIn , \s14.dbus_out , \s14.en , \s14.Tdone  );
  input [63:0] \m0.addrM64 ;
  input [63:0] \m0.DoutM ;
  output [63:0] \m0.MinData ;
  output [63:0] \s0.addr ;
  output [63:0] \s0.SbusIn ;
  input [63:0] \s0.dbus_out ;
  input [63:0] \m1.addrM64 ;
  input [63:0] \m1.DoutM ;
  output [63:0] \m1.MinData ;
  output [63:0] \s1.addr ;
  output [63:0] \s1.SbusIn ;
  input [63:0] \s1.dbus_out ;
  input [63:0] \m2.addrM64 ;
  input [63:0] \m2.DoutM ;
  output [63:0] \m2.MinData ;
  output [63:0] \s2.addr ;
  output [63:0] \s2.SbusIn ;
  input [63:0] \s2.dbus_out ;
  input [63:0] \m3.addrM64 ;
  input [63:0] \m3.DoutM ;
  output [63:0] \m3.MinData ;
  output [63:0] \s3.addr ;
  output [63:0] \s3.SbusIn ;
  input [63:0] \s3.dbus_out ;
  input [63:0] \m4.addrM64 ;
  input [63:0] \m4.DoutM ;
  output [63:0] \m4.MinData ;
  output [63:0] \s4.addr ;
  output [63:0] \s4.SbusIn ;
  input [63:0] \s4.dbus_out ;
  input [63:0] \m5.addrM64 ;
  input [63:0] \m5.DoutM ;
  output [63:0] \m5.MinData ;
  output [63:0] \s5.addr ;
  output [63:0] \s5.SbusIn ;
  input [63:0] \s5.dbus_out ;
  input [63:0] \m6.addrM64 ;
  input [63:0] \m6.DoutM ;
  output [63:0] \m6.MinData ;
  output [63:0] \s6.addr ;
  output [63:0] \s6.SbusIn ;
  input [63:0] \s6.dbus_out ;
  output [63:0] \s7.addr ;
  output [63:0] \s7.SbusIn ;
  input [63:0] \s7.dbus_out ;
  output [63:0] \s8.addr ;
  output [63:0] \s8.SbusIn ;
  input [63:0] \s8.dbus_out ;
  output [63:0] \s9.addr ;
  output [63:0] \s9.SbusIn ;
  input [63:0] \s9.dbus_out ;
  output [63:0] \s10.addr ;
  output [63:0] \s10.SbusIn ;
  input [63:0] \s10.dbus_out ;
  output [63:0] \s11.addr ;
  output [63:0] \s11.SbusIn ;
  input [63:0] \s11.dbus_out ;
  output [63:0] \s12.addr ;
  output [63:0] \s12.SbusIn ;
  input [63:0] \s12.dbus_out ;
  output [63:0] \s13.addr ;
  output [63:0] \s13.SbusIn ;
  input [63:0] \s13.dbus_out ;
  output [63:0] \s14.addr ;
  output [63:0] \s14.SbusIn ;
  input [63:0] \s14.dbus_out ;
  input \c1.sysClk , \c1.Breset , \m0.need , \m1.need , \m2.need , \m3.need ,
         \m4.need , \m5.need , \m6.need ;
  output \m0.ack , \m0.Tdone_mstr , \s0.en , \s0.Tdone , \m1.ack ,
         \m1.Tdone_mstr , \s1.en , \s1.Tdone , \m2.ack , \m2.Tdone_mstr ,
         \s2.en , \s2.Tdone , \m3.ack , \m3.Tdone_mstr , \s3.en , \s3.Tdone ,
         \m4.ack , \m4.Tdone_mstr , \s4.en , \s4.Tdone , \m5.ack ,
         \m5.Tdone_mstr , \s5.en , \s5.Tdone , \m6.ack , \m6.Tdone_mstr ,
         \s6.en , \s6.Tdone , \s7.en , \s7.Tdone , \s8.en , \s8.Tdone ,
         \s9.en , \s9.Tdone , \s10.en , \s10.Tdone , \s11.en , \s11.Tdone ,
         \s12.en , \s12.Tdone , \s13.en , \s13.Tdone , \s14.en , \s14.Tdone ;
  wire   \nx_st[2] , n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, \s13.addr[13] , n3405, n3406, n3407,
         n3408, n3409, n3410, \s13.addr[18] , n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, \s8.addr[17] , n4386, \s4.en ,
         \s4.addr[14] , \s8.addr[15] , \s8.en , \s12.addr[10] , \s3.addr[9] ,
         \s3.addr[14] , \s11.addr[19] , \s7.addr[19] , \s7.en , \s12.addr[11] ,
         \s5.addr[14] , \s9.addr[8] , \s6.en , n4405, \s2.addr[19] ,
         \s9.addr[7] , \s2.addr[16] , \s11.addr[17] , \s10.en , \s14.addr[18] ,
         \s10.addr[9] , n4418, n4419, n4420, n4421, n4422, \s14.addr[16] ,
         \s1.addr[17] , \s1.en , \s1.addr[15] , \s12.addr[16] , \s13.addr[15] ,
         \s0.addr[17] , n5445, n5518, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, \s9.addr[16] ,
         n5590, \s7.addr[16] , \s14.addr[17] ;
  wire   [63:0] data_stm_d;
  assign \s0.addr  [16] = 1'b0;
  assign \s0.addr  [11] = 1'b0;
  assign \s0.addr  [7] = 1'b0;
  assign \s1.addr  [10] = 1'b0;
  assign \s2.addr  [15] = 1'b0;
  assign \s2.addr  [14] = 1'b0;
  assign \s3.addr  [15] = 1'b0;
  assign \s3.addr  [10] = 1'b0;
  assign \s4.addr  [10] = 1'b0;
  assign \s6.addr  [14] = 1'b0;
  assign \s6.addr  [9] = 1'b0;
  assign \s6.addr  [7] = 1'b0;
  assign \s8.addr  [13] = 1'b0;
  assign \s8.addr  [10] = 1'b0;
  assign \s9.addr  [14] = 1'b0;
  assign \s9.addr  [9] = 1'b0;
  assign \s10.addr  [14] = 1'b0;
  assign \s10.addr  [10] = 1'b0;
  assign \s0.addr  [15] = 1'b0;
  assign \s0.addr  [8] = 1'b0;
  assign \s4.addr  [16] = 1'b0;
  assign \s4.addr  [8] = 1'b0;
  assign \s5.addr  [11] = 1'b0;
  assign \s5.addr  [9] = 1'b0;
  assign \s5.addr  [8] = 1'b0;
  assign \s6.addr  [16] = 1'b0;
  assign \s6.addr  [12] = 1'b0;
  assign \s14.addr  [15] = 1'b0;
  assign \s14.addr  [12] = 1'b0;
  assign \s1.addr  [13] = 1'b0;
  assign \s1.addr  [11] = 1'b0;
  assign \s2.addr  [13] = 1'b0;
  assign \s2.addr  [11] = 1'b0;
  assign \s2.addr  [10] = 1'b0;
  assign \s2.addr  [9] = 1'b0;
  assign \s3.addr  [13] = 1'b0;
  assign \s3.addr  [12] = 1'b0;
  assign \s3.addr  [11] = 1'b0;
  assign \s4.addr  [11] = 1'b0;
  assign \s5.addr  [16] = 1'b0;
  assign \s5.addr  [15] = 1'b0;
  assign \s7.addr  [15] = 1'b0;
  assign \s7.addr  [14] = 1'b0;
  assign \s9.addr  [12] = 1'b0;
  assign \s10.addr  [12] = 1'b0;
  assign \s10.addr  [11] = 1'b0;
  assign \s12.addr  [15] = 1'b0;
  assign \s12.addr  [13] = 1'b0;
  assign \s13.addr  [14] = 1'b0;
  assign \s14.addr  [13] = 1'b0;
  assign \s14.addr  [10] = 1'b0;
  assign \s13.en  = \s13.addr[13] ;
  assign \s13.addr  [13] = \s13.addr[13] ;
  assign \s13.addr  [17] = \s13.addr[18] ;
  assign \s13.addr  [18] = \s13.addr[18] ;
  assign \s8.addr  [16] = \s8.addr[17] ;
  assign \s8.addr  [17] = \s8.addr[17] ;
  assign \s4.addr  [17] = \s4.en ;
  assign \s4.addr  [12] = \s4.en ;
  assign \s4.addr  [9] = \s4.en ;
  assign \s4.addr  [15] = \s4.addr[14] ;
  assign \s4.addr  [13] = \s4.addr[14] ;
  assign \s4.addr  [18] = \s4.addr[14] ;
  assign \s4.addr  [14] = \s4.addr[14] ;
  assign \s8.addr  [12] = \s8.addr[15] ;
  assign \s8.addr  [14] = \s8.addr[15] ;
  assign \s8.addr  [15] = \s8.addr[15] ;
  assign \s8.addr  [11] = \s8.en ;
  assign \s8.addr  [19] = \s8.en ;
  assign \s8.addr  [18] = \s8.en ;
  assign \s12.addr  [9] = \s12.addr[10] ;
  assign \s12.addr  [14] = \s12.addr[10] ;
  assign \s12.addr  [10] = \s12.addr[10] ;
  assign \s3.addr  [17] = \s3.addr[9] ;
  assign \s3.addr  [9] = \s3.addr[9] ;
  assign \s3.en  = \s3.addr[14] ;
  assign \s3.addr  [16] = \s3.addr[14] ;
  assign \s3.addr  [19] = \s3.addr[14] ;
  assign \s3.addr  [14] = \s3.addr[14] ;
  assign \s11.addr  [13] = \s11.addr[19] ;
  assign \s11.addr  [12] = \s11.addr[19] ;
  assign \s11.addr  [15] = \s11.addr[19] ;
  assign \s11.addr  [19] = \s11.addr[19] ;
  assign \s7.addr  [12] = \s7.addr[19] ;
  assign \s7.addr  [19] = \s7.addr[19] ;
  assign \s7.addr  [17] = \s7.en ;
  assign \s7.addr  [18] = \s7.en ;
  assign \s12.addr  [12] = \s12.addr[11] ;
  assign \s12.addr  [11] = \s12.addr[11] ;
  assign \s5.en  = \s5.addr[14] ;
  assign \s5.addr  [10] = \s5.addr[14] ;
  assign \s5.addr  [19] = \s5.addr[14] ;
  assign \s5.addr  [18] = \s5.addr[14] ;
  assign \s5.addr  [17] = \s5.addr[14] ;
  assign \s5.addr  [12] = \s5.addr[14] ;
  assign \s5.addr  [13] = \s5.addr[14] ;
  assign \s5.addr  [14] = \s5.addr[14] ;
  assign \s9.addr  [10] = \s9.addr[8] ;
  assign \s9.addr  [13] = \s9.addr[8] ;
  assign \s9.addr  [17] = \s9.addr[8] ;
  assign \s9.addr  [8] = \s9.addr[8] ;
  assign \s6.addr  [11] = \s6.en ;
  assign \s6.addr  [8] = \s6.en ;
  assign \s6.addr  [13] = \s6.en ;
  assign \s6.addr  [18] = \s6.en ;
  assign \s6.addr  [15] = \s6.en ;
  assign \s6.addr  [10] = \s6.en ;
  assign \s6.addr  [19] = \s6.en ;
  assign \s2.addr  [12] = \s2.addr[19] ;
  assign \s2.addr  [19] = \s2.addr[19] ;
  assign \s9.addr  [11] = \s9.addr[7] ;
  assign \s9.addr  [7] = \s9.addr[7] ;
  assign \s2.en  = \s2.addr[16] ;
  assign \s2.addr  [18] = \s2.addr[16] ;
  assign \s2.addr  [17] = \s2.addr[16] ;
  assign \s2.addr  [16] = \s2.addr[16] ;
  assign \s11.addr  [16] = \s11.addr[17] ;
  assign \s11.addr  [14] = \s11.addr[17] ;
  assign \s11.addr  [18] = \s11.addr[17] ;
  assign \s11.addr  [17] = \s11.addr[17] ;
  assign \s10.addr  [16] = \s10.en ;
  assign \s10.addr  [15] = \s10.en ;
  assign \s10.addr  [18] = \s10.en ;
  assign \s10.addr  [13] = \s10.en ;
  assign \s14.addr  [9] = \s14.addr[18] ;
  assign \s14.en  = \s14.addr[18] ;
  assign \s14.addr  [18] = \s14.addr[18] ;
  assign \s10.addr  [19] = \s10.addr[9] ;
  assign \s10.addr  [9] = \s10.addr[9] ;
  assign \s14.addr  [14] = \s14.addr[16] ;
  assign \s14.addr  [16] = \s14.addr[16] ;
  assign \s1.addr  [9] = \s1.addr[17] ;
  assign \s1.addr  [18] = \s1.addr[17] ;
  assign \s1.addr  [14] = \s1.addr[17] ;
  assign \s1.addr  [17] = \s1.addr[17] ;
  assign \s1.addr  [8] = \s1.en ;
  assign \s1.addr  [16] = \s1.addr[15] ;
  assign \s1.addr  [12] = \s1.addr[15] ;
  assign \s1.addr  [15] = \s1.addr[15] ;
  assign \s12.addr  [18] = \s12.addr[16] ;
  assign \s12.addr  [17] = \s12.addr[16] ;
  assign \s12.en  = \s12.addr[16] ;
  assign \s12.addr  [16] = \s12.addr[16] ;
  assign \s13.addr  [16] = \s13.addr[15] ;
  assign \s13.addr  [19] = \s13.addr[15] ;
  assign \s13.addr  [12] = \s13.addr[15] ;
  assign \s13.addr  [15] = \s13.addr[15] ;
  assign \s0.addr  [19] = \s0.addr[17] ;
  assign \s0.addr  [18] = \s0.addr[17] ;
  assign \s0.addr  [10] = \s0.addr[17] ;
  assign \s0.addr  [9] = \s0.addr[17] ;
  assign \s0.addr  [17] = \s0.addr[17] ;
  assign \s9.addr  [19] = \s9.addr[16] ;
  assign \s9.addr  [18] = \s9.addr[16] ;
  assign \s9.addr  [16] = \s9.addr[16] ;
  assign \s7.addr  [13] = \s7.addr[16] ;
  assign \s7.addr  [16] = \s7.addr[16] ;
  assign \s14.addr  [19] = \s14.addr[17] ;
  assign \s14.addr  [17] = \s14.addr[17] ;

  CFDN4QX4 \st_reg[0]  ( .D(n4421), .CPN(\c1.sysClk ), .SD(n5518), .Q(n4422)
         );
  CFDN4QX4 \st_reg[2]  ( .D(\nx_st[2] ), .CPN(\c1.sysClk ), .SD(n5518), .Q(
        n4420) );
  CFDN4QX4 \st_reg[1]  ( .D(n4418), .CPN(\c1.sysClk ), .SD(n5518), .Q(n4419)
         );
  CFDN1XL \data_stm_d_reg[17]  ( .D(n1737), .CPN(\c1.sysClk ), .Q(
        data_stm_d[17]), .QN(n5540) );
  CFDN1XL \data_stm_d_reg[62]  ( .D(n1692), .CPN(n4386), .Q(data_stm_d[62]), 
        .QN(n5586) );
  CFDN1XL \data_stm_d_reg[33]  ( .D(n1721), .CPN(n4386), .Q(data_stm_d[33]), 
        .QN(n5556) );
  CFDN1XL \data_stm_d_reg[59]  ( .D(n1695), .CPN(n4386), .Q(data_stm_d[59]), 
        .QN(n5583) );
  CFDN1XL \data_stm_d_reg[58]  ( .D(n1696), .CPN(n4386), .Q(data_stm_d[58]), 
        .QN(n5582) );
  CFDN1XL \data_stm_d_reg[50]  ( .D(n1704), .CPN(n4386), .Q(data_stm_d[50]), 
        .QN(n5574) );
  CFDN1XL \data_stm_d_reg[19]  ( .D(n1735), .CPN(n4386), .Q(data_stm_d[19]), 
        .QN(n5542) );
  CFDN1XL \data_stm_d_reg[37]  ( .D(n1717), .CPN(n4386), .Q(data_stm_d[37]), 
        .QN(n5560) );
  CFDN1XL \data_stm_d_reg[28]  ( .D(n1726), .CPN(n4386), .Q(data_stm_d[28]), 
        .QN(n5551) );
  CFDN1XL \data_stm_d_reg[25]  ( .D(n1729), .CPN(n4386), .Q(data_stm_d[25]), 
        .QN(n5548) );
  CFDN1XL \data_stm_d_reg[32]  ( .D(n1722), .CPN(n4386), .Q(data_stm_d[32]), 
        .QN(n5555) );
  CFDN1XL \data_stm_d_reg[27]  ( .D(n1727), .CPN(n4386), .Q(data_stm_d[27]), 
        .QN(n5550) );
  CFDN1XL \data_stm_d_reg[16]  ( .D(n1738), .CPN(n4386), .Q(data_stm_d[16]), 
        .QN(n5539) );
  CFDN1XL \data_stm_d_reg[63]  ( .D(n1691), .CPN(n4386), .Q(data_stm_d[63]), 
        .QN(n5587) );
  CFDN1XL \data_stm_d_reg[42]  ( .D(n1712), .CPN(n4386), .Q(data_stm_d[42]), 
        .QN(n5565) );
  CFDN1XL \data_stm_d_reg[30]  ( .D(n1724), .CPN(n4386), .Q(data_stm_d[30]), 
        .QN(n5553) );
  CFDN1XL \data_stm_d_reg[24]  ( .D(n1730), .CPN(n4386), .Q(data_stm_d[24]), 
        .QN(n5547) );
  CFDN1XL \data_stm_d_reg[53]  ( .D(n1701), .CPN(n4386), .Q(data_stm_d[53]), 
        .QN(n5577) );
  CFDN1XL \data_stm_d_reg[36]  ( .D(n1718), .CPN(n4386), .Q(data_stm_d[36]), 
        .QN(n5559) );
  CFDN1XL \data_stm_d_reg[39]  ( .D(n1715), .CPN(n4386), .Q(data_stm_d[39]), 
        .QN(n5562) );
  CFDN1XL \data_stm_d_reg[31]  ( .D(n1723), .CPN(n4386), .Q(data_stm_d[31]), 
        .QN(n5554) );
  CFDN1XL \data_stm_d_reg[34]  ( .D(n1720), .CPN(n4386), .Q(data_stm_d[34]), 
        .QN(n5557) );
  CFDN1XL \data_stm_d_reg[56]  ( .D(n1698), .CPN(n4386), .Q(data_stm_d[56]), 
        .QN(n5580) );
  CFDN1XL \data_stm_d_reg[48]  ( .D(n1706), .CPN(n4386), .Q(data_stm_d[48]), 
        .QN(n5571) );
  CFDN1XL \data_stm_d_reg[20]  ( .D(n1734), .CPN(n4386), .Q(data_stm_d[20]), 
        .QN(n5543) );
  CFDN1XL \data_stm_d_reg[12]  ( .D(n1742), .CPN(\c1.sysClk ), .Q(
        data_stm_d[12]), .QN(n5535) );
  CFDN1XL \data_stm_d_reg[1]  ( .D(n1753), .CPN(\c1.sysClk ), .Q(data_stm_d[1]), .QN(n5524) );
  CFDN1XL \data_stm_d_reg[6]  ( .D(n1748), .CPN(\c1.sysClk ), .Q(data_stm_d[6]), .QN(n5529) );
  CFDN1XL \data_stm_d_reg[10]  ( .D(n1744), .CPN(\c1.sysClk ), .Q(
        data_stm_d[10]), .QN(n5533) );
  CFDN1XL \data_stm_d_reg[13]  ( .D(n1741), .CPN(\c1.sysClk ), .Q(
        data_stm_d[13]), .QN(n5536) );
  CFDN1XL \data_stm_d_reg[8]  ( .D(n1746), .CPN(\c1.sysClk ), .Q(data_stm_d[8]), .QN(n5531) );
  CFDN1XL \data_stm_d_reg[0]  ( .D(n1754), .CPN(\c1.sysClk ), .Q(data_stm_d[0]), .QN(n5523) );
  CFDN1XL \data_stm_d_reg[15]  ( .D(n1739), .CPN(\c1.sysClk ), .Q(
        data_stm_d[15]), .QN(n5538) );
  CFDN1XL \data_stm_d_reg[61]  ( .D(n1693), .CPN(n4386), .Q(data_stm_d[61]), 
        .QN(n5585) );
  CFDN1XL \data_stm_d_reg[47]  ( .D(n1707), .CPN(n4386), .Q(data_stm_d[47]), 
        .QN(n5570) );
  CFDN1XL \data_stm_d_reg[45]  ( .D(n1709), .CPN(n4386), .Q(data_stm_d[45]), 
        .QN(n5568) );
  CFDN1XL \data_stm_d_reg[44]  ( .D(n1710), .CPN(n4386), .Q(data_stm_d[44]), 
        .QN(n5567) );
  CFDN1XL \data_stm_d_reg[41]  ( .D(n1713), .CPN(n4386), .Q(data_stm_d[41]), 
        .QN(n5564) );
  CFDN1XL \data_stm_d_reg[40]  ( .D(n1714), .CPN(n4386), .Q(data_stm_d[40]), 
        .QN(n5563) );
  CFDN1XL \data_stm_d_reg[60]  ( .D(n1694), .CPN(n4386), .Q(data_stm_d[60]), 
        .QN(n5584) );
  CFDN1XL \data_stm_d_reg[57]  ( .D(n1697), .CPN(n4386), .Q(data_stm_d[57]), 
        .QN(n5581) );
  CFDN1XL \data_stm_d_reg[55]  ( .D(n1699), .CPN(n4386), .Q(data_stm_d[55]), 
        .QN(n5579) );
  CFDN1XL \data_stm_d_reg[54]  ( .D(n1700), .CPN(n4386), .Q(data_stm_d[54]), 
        .QN(n5578) );
  CFDN1XL \data_stm_d_reg[52]  ( .D(n1702), .CPN(n4386), .Q(data_stm_d[52]), 
        .QN(n5576) );
  CFDN1XL \data_stm_d_reg[51]  ( .D(n1703), .CPN(n4386), .Q(data_stm_d[51]), 
        .QN(n5575) );
  CFDN1XL \data_stm_d_reg[49]  ( .D(n1705), .CPN(n4386), .Q(data_stm_d[49]), 
        .QN(n5572) );
  CFDN1XL \data_stm_d_reg[46]  ( .D(n1708), .CPN(n4386), .Q(data_stm_d[46]), 
        .QN(n5569) );
  CFDN1XL \data_stm_d_reg[43]  ( .D(n1711), .CPN(n4386), .Q(data_stm_d[43]), 
        .QN(n5566) );
  CFDN1XL \data_stm_d_reg[38]  ( .D(n1716), .CPN(n4386), .Q(data_stm_d[38]), 
        .QN(n5561) );
  CFDN1XL \data_stm_d_reg[35]  ( .D(n1719), .CPN(n4386), .Q(data_stm_d[35]), 
        .QN(n5558) );
  CFDN1XL \data_stm_d_reg[29]  ( .D(n1725), .CPN(n4386), .Q(data_stm_d[29]), 
        .QN(n5552) );
  CFDN1XL \data_stm_d_reg[26]  ( .D(n1728), .CPN(n4386), .Q(data_stm_d[26]), 
        .QN(n5549) );
  CFDN1XL \data_stm_d_reg[23]  ( .D(n1731), .CPN(n4386), .Q(data_stm_d[23]), 
        .QN(n5546) );
  CFDN1XL \data_stm_d_reg[22]  ( .D(n1732), .CPN(n4386), .Q(data_stm_d[22]), 
        .QN(n5545) );
  CFDN1XL \data_stm_d_reg[21]  ( .D(n1733), .CPN(n4386), .Q(data_stm_d[21]), 
        .QN(n5544) );
  CFDN1XL \data_stm_d_reg[18]  ( .D(n1736), .CPN(n4386), .Q(data_stm_d[18]), 
        .QN(n5541) );
  CFDN1XL \data_stm_d_reg[7]  ( .D(n1747), .CPN(\c1.sysClk ), .Q(data_stm_d[7]), .QN(n5530) );
  CFDN1XL \data_stm_d_reg[5]  ( .D(n1749), .CPN(\c1.sysClk ), .Q(data_stm_d[5]), .QN(n5528) );
  CFDN1XL \data_stm_d_reg[4]  ( .D(n1750), .CPN(\c1.sysClk ), .Q(data_stm_d[4]), .QN(n5527) );
  CFDN1XL \data_stm_d_reg[3]  ( .D(n1751), .CPN(\c1.sysClk ), .Q(data_stm_d[3]), .QN(n5526) );
  CFDN1XL \data_stm_d_reg[2]  ( .D(n1752), .CPN(\c1.sysClk ), .Q(data_stm_d[2]), .QN(n5525) );
  CFDN1XL \data_stm_d_reg[14]  ( .D(n1740), .CPN(\c1.sysClk ), .Q(
        data_stm_d[14]), .QN(n5537) );
  CFDN1XL \data_stm_d_reg[11]  ( .D(n1743), .CPN(\c1.sysClk ), .Q(
        data_stm_d[11]), .QN(n5534) );
  CFDN1XL \data_stm_d_reg[9]  ( .D(n1745), .CPN(\c1.sysClk ), .Q(data_stm_d[9]), .QN(n5532) );
  CND2X1 U4138 ( .A(n1997), .B(n1992), .Z(n1890) );
  CND2X2 U4139 ( .A(n1933), .B(\m0.addrM64 [3]), .Z(n1993) );
  CIVX2 U4140 ( .A(n2780), .Z(n2788) );
  COND1X2 U4141 ( .A(n3476), .B(n1980), .C(n3409), .Z(n1981) );
  CND3X2 U4142 ( .A(n2465), .B(n2783), .C(n2093), .Z(n2129) );
  CND2IX2 U4143 ( .B(n3478), .A(n2623), .Z(n2522) );
  CND3X1 U4144 ( .A(n3454), .B(n2728), .C(n5518), .Z(n2734) );
  CND2X1 U4145 ( .A(n1904), .B(\m5.addrM64 [2]), .Z(n2632) );
  CND2X1 U4146 ( .A(n2252), .B(\m4.addrM64 [1]), .Z(n1908) );
  CND2X2 U4147 ( .A(n1977), .B(n1976), .Z(n2116) );
  CNR2X1 U4148 ( .A(n2188), .B(n2187), .Z(n2190) );
  CND2X1 U4149 ( .A(n2246), .B(\m6.addrM64 [18]), .Z(n2048) );
  CNR2IX1 U4150 ( .B(\m5.addrM64 [19]), .A(n2248), .Z(n2036) );
  CAN2X1 U4151 ( .A(n2774), .B(n2773), .Z(n2777) );
  CNR2X1 U4152 ( .A(n2613), .B(\c1.Breset ), .Z(n2615) );
  CNR2IX1 U4153 ( .B(n2762), .A(n3405), .Z(n2461) );
  CAN2X1 U4154 ( .A(n2780), .B(n4326), .Z(n2642) );
  CND2X2 U4155 ( .A(n2217), .B(n2783), .Z(n2218) );
  CND2X1 U4156 ( .A(n2088), .B(\m1.addrM64 [6]), .Z(n1942) );
  CND2X2 U4157 ( .A(n2089), .B(\m5.addrM64 [4]), .Z(n2002) );
  CND2X2 U4158 ( .A(n2089), .B(\m5.addrM64 [8]), .Z(n1879) );
  CNR2X1 U4159 ( .A(n2050), .B(n2049), .Z(n2052) );
  CNR2IX1 U4160 ( .B(\m4.addrM64 [18]), .A(n2078), .Z(n2049) );
  CND2X1 U4161 ( .A(n2048), .B(n2047), .Z(n2050) );
  CANR2X1 U4162 ( .A(n2245), .B(\m0.addrM64 [17]), .C(\m5.addrM64 [17]), .D(
        n2089), .Z(n2041) );
  CND2X1 U4163 ( .A(n2088), .B(\m1.addrM64 [12]), .Z(n2075) );
  CND3X2 U4164 ( .A(n1988), .B(n1984), .C(n1987), .Z(n2198) );
  CND2X2 U4165 ( .A(n2252), .B(\m4.addrM64 [4]), .Z(n2108) );
  CANR2X1 U4166 ( .A(n2085), .B(\m2.addrM64 [12]), .C(\m6.addrM64 [12]), .D(
        n2246), .Z(n2081) );
  CND3X2 U4167 ( .A(n1875), .B(n1874), .C(n1873), .Z(n2201) );
  CND3X1 U4168 ( .A(n2793), .B(n2788), .C(n2125), .Z(n2127) );
  COR2X1 U4169 ( .A(n2761), .B(n2031), .Z(n2094) );
  CND2X1 U4170 ( .A(n2180), .B(n2623), .Z(n2182) );
  CND2X2 U4171 ( .A(n2458), .B(n2457), .Z(n2512) );
  COND1X1 U4172 ( .A(n2456), .B(n2522), .C(n4257), .Z(n2458) );
  CND2X1 U4173 ( .A(n2547), .B(n2545), .Z(n2525) );
  COR2X1 U4174 ( .A(n2736), .B(n2735), .Z(n2737) );
  CNR3X2 U4175 ( .A(n2734), .B(n2733), .C(n2732), .Z(n2738) );
  CND2X2 U4176 ( .A(n2001), .B(n2000), .Z(n2772) );
  CNR2X1 U4177 ( .A(n1999), .B(n1998), .Z(n2000) );
  CND2IX1 U4178 ( .B(n2757), .A(n2756), .Z(n2758) );
  CND3XL U4179 ( .A(n2753), .B(n2752), .C(n2751), .Z(n2759) );
  CND2X2 U4180 ( .A(n1934), .B(n1973), .Z(n1935) );
  CND2X1 U4181 ( .A(n2855), .B(\m3.addrM64 [6]), .Z(n1948) );
  CND2X2 U4182 ( .A(n2088), .B(\m1.addrM64 [4]), .Z(n2111) );
  CIVDX1 U4183 ( .A(n2108), .Z0(n1959), .Z1(n2110) );
  CND2X1 U4184 ( .A(n2246), .B(\m6.addrM64 [8]), .Z(n1883) );
  CND2X1 U4185 ( .A(n2088), .B(\m1.addrM64 [8]), .Z(n1884) );
  CND2X1 U4186 ( .A(n1961), .B(\m6.addrM64 [10]), .Z(n1862) );
  CND2X1 U4187 ( .A(\m1.addrM64 [16]), .B(n2088), .Z(n2068) );
  CNIVX1 U4188 ( .A(\s3.addr[14] ), .Z(n4101) );
  CIVX2 U4189 ( .A(n2116), .Z(n1978) );
  CIVX2 U4190 ( .A(n2117), .Z(n1979) );
  CIVX2 U4191 ( .A(n3448), .Z(n3484) );
  CND2X2 U4192 ( .A(n2196), .B(n2195), .Z(n2452) );
  CIVX2 U4193 ( .A(\m5.ack ), .Z(n2979) );
  CND3X1 U4194 ( .A(n2282), .B(n2281), .C(n2280), .Z(n4200) );
  CANR1XL U4195 ( .A(n3434), .B(\m0.DoutM [3]), .C(n2279), .Z(n2280) );
  COND1XL U4196 ( .A(n3432), .B(n3060), .C(n3059), .Z(n3064) );
  CANR1XL U4197 ( .A(\m0.DoutM [7]), .B(n3434), .C(n2438), .Z(n2439) );
  CANR1XL U4198 ( .A(n3431), .B(\m1.DoutM [7]), .C(n2436), .Z(n2442) );
  CANR1XL U4199 ( .A(n3431), .B(\m1.DoutM [16]), .C(n3260), .Z(n3265) );
  COND1XL U4200 ( .A(n3432), .B(n2347), .C(n2346), .Z(n2351) );
  COND1XL U4201 ( .A(n2349), .B(n3439), .C(n2348), .Z(n2350) );
  CANR1XL U4202 ( .A(n3431), .B(\m1.DoutM [21]), .C(n2980), .Z(n2985) );
  CANR1XL U4203 ( .A(n3434), .B(\m0.DoutM [24]), .C(n2952), .Z(n2958) );
  COND1XL U4204 ( .A(n3432), .B(n2366), .C(n2365), .Z(n2370) );
  COND1XL U4205 ( .A(n2368), .B(n3439), .C(n2367), .Z(n2369) );
  CANR1XL U4206 ( .A(n3431), .B(\m1.DoutM [26]), .C(n2556), .Z(n2561) );
  COND1XL U4207 ( .A(n3432), .B(n2871), .C(n2870), .Z(n2873) );
  CND3X1 U4208 ( .A(n2885), .B(n2884), .C(n2883), .Z(n4197) );
  COND1XL U4209 ( .A(n3432), .B(n2879), .C(n2878), .Z(n2880) );
  CND3X1 U4210 ( .A(n2396), .B(n2395), .C(n2394), .Z(n4145) );
  COND1XL U4211 ( .A(n3432), .B(n2390), .C(n2389), .Z(n2391) );
  COND1XL U4212 ( .A(n3432), .B(n3079), .C(n3078), .Z(n3081) );
  CND3X1 U4213 ( .A(n2601), .B(n2600), .C(n2599), .Z(n4171) );
  COND1XL U4214 ( .A(n3432), .B(n2595), .C(n2594), .Z(n2596) );
  CND3X1 U4215 ( .A(n2611), .B(n2610), .C(n2609), .Z(n4178) );
  COND1XL U4216 ( .A(n3432), .B(n2605), .C(n2604), .Z(n2606) );
  CANR1XL U4217 ( .A(n3434), .B(\m0.DoutM [36]), .C(n2988), .Z(n2989) );
  COND1XL U4218 ( .A(n3432), .B(n3233), .C(n3232), .Z(n3234) );
  CANR1XL U4219 ( .A(n3434), .B(\m0.DoutM [43]), .C(n3227), .Z(n3228) );
  CANR1XL U4220 ( .A(n3434), .B(\m0.DoutM [44]), .C(n2518), .Z(n2519) );
  COND1XL U4221 ( .A(n3432), .B(n3323), .C(n3322), .Z(n3327) );
  COND1XL U4222 ( .A(n3325), .B(n3439), .C(n3324), .Z(n3326) );
  CANR1XL U4223 ( .A(n3434), .B(\m0.DoutM [46]), .C(n2415), .Z(n2416) );
  CANR1XL U4224 ( .A(n3434), .B(\m0.DoutM [53]), .C(n2423), .Z(n2424) );
  CND3X1 U4225 ( .A(n3349), .B(n3348), .C(n3347), .Z(n4159) );
  COND1XL U4226 ( .A(n3432), .B(n3343), .C(n3342), .Z(n3344) );
  CANR1XL U4227 ( .A(n3431), .B(\m1.DoutM [57]), .C(n3358), .Z(n3365) );
  CANR1XL U4228 ( .A(\m3.DoutM [57]), .B(n3361), .C(n3360), .Z(n3363) );
  CANR1XL U4229 ( .A(n3434), .B(\m0.DoutM [58]), .C(n3197), .Z(n3201) );
  CANR1XL U4230 ( .A(\m1.DoutM [58]), .B(n3431), .C(n3196), .Z(n3202) );
  CANR1XL U4231 ( .A(n3434), .B(\m0.DoutM [59]), .C(n2499), .Z(n2500) );
  COND1XL U4232 ( .A(n3432), .B(n2678), .C(n2677), .Z(n2680) );
  CANR1XL U4233 ( .A(n3434), .B(\m0.DoutM [63]), .C(n3215), .Z(n3221) );
  CNR2X1 U4234 ( .A(n2635), .B(n2634), .Z(n2636) );
  CAN2X1 U4235 ( .A(n2633), .B(n2632), .Z(n2638) );
  CANR1XL U4236 ( .A(n3434), .B(\m0.addrM64 [21]), .C(n2566), .Z(n2567) );
  CANR1XL U4237 ( .A(n3431), .B(\m1.addrM64 [22]), .C(n3276), .Z(n3281) );
  CND3X1 U4238 ( .A(n3141), .B(n3140), .C(n3139), .Z(n4118) );
  COND1XL U4239 ( .A(n3432), .B(n3134), .C(n3133), .Z(n3135) );
  CND3X1 U4240 ( .A(n3250), .B(n3249), .C(n3248), .Z(n4199) );
  COND1XL U4241 ( .A(n3432), .B(n3244), .C(n3243), .Z(n3245) );
  COND1XL U4242 ( .A(n3432), .B(n2909), .C(n2908), .Z(n2913) );
  COND1XL U4243 ( .A(n2911), .B(n3439), .C(n2910), .Z(n2912) );
  CANR1XL U4244 ( .A(n3431), .B(\m1.addrM64 [36]), .C(n2706), .Z(n2711) );
  CND3X1 U4245 ( .A(n3094), .B(n3093), .C(n3092), .Z(n4177) );
  COND1XL U4246 ( .A(n3432), .B(n3087), .C(n3086), .Z(n3088) );
  CND2X1 U4247 ( .A(n3310), .B(n3309), .Z(n3486) );
  COND1XL U4248 ( .A(n3432), .B(n3304), .C(n3303), .Z(n3308) );
  CANR1XL U4249 ( .A(n3434), .B(\m0.addrM64 [42]), .C(n3172), .Z(n3178) );
  COND1XL U4250 ( .A(n3432), .B(n2844), .C(n2843), .Z(n2848) );
  CANR1XL U4251 ( .A(\m0.addrM64 [46]), .B(n3434), .C(n2835), .Z(n2836) );
  CANR1XL U4252 ( .A(n3431), .B(\m1.addrM64 [46]), .C(n2833), .Z(n2839) );
  CND3X1 U4253 ( .A(n2969), .B(n2968), .C(n2967), .Z(n4155) );
  COND1XL U4254 ( .A(n3432), .B(n2963), .C(n2962), .Z(n2964) );
  CND3X1 U4255 ( .A(n3130), .B(n3129), .C(n3128), .Z(n4164) );
  COND1XL U4256 ( .A(n3432), .B(n3124), .C(n3123), .Z(n3125) );
  CANR1XL U4257 ( .A(\m1.addrM64 [52]), .B(n3431), .C(n3180), .Z(n3187) );
  CND3X1 U4258 ( .A(n3275), .B(n3274), .C(n3273), .Z(n4174) );
  CANR1XL U4259 ( .A(n3431), .B(\m1.addrM64 [53]), .C(n3272), .Z(n3274) );
  CND2X1 U4260 ( .A(n3371), .B(\m3.addrM64 [53]), .Z(n3273) );
  COND1XL U4261 ( .A(n3432), .B(n3269), .C(n3268), .Z(n3270) );
  COND1XL U4262 ( .A(n3432), .B(n2667), .C(n2666), .Z(n2671) );
  COND1XL U4263 ( .A(n2669), .B(n3439), .C(n2668), .Z(n2670) );
  CANR1XL U4264 ( .A(n3431), .B(\m1.addrM64 [56]), .C(n2658), .Z(n2662) );
  CND3X1 U4265 ( .A(n2946), .B(n2945), .C(n2944), .Z(n3477) );
  CANR1XL U4266 ( .A(n3431), .B(\m1.addrM64 [62]), .C(n2947), .Z(n2951) );
  CANR1XL U4267 ( .A(\m1.addrM64 [63]), .B(n3431), .C(n3421), .Z(n3429) );
  CIVX3 U4268 ( .A(\m1.ack ), .Z(n3383) );
  CNIVX8 U4269 ( .A(n2247), .Z(n3431) );
  CIVDX1 U4270 ( .A(n4338), .Z0(n4254), .Z1(n4334) );
  CIVX2 U4271 ( .A(n2199), .Z(n4335) );
  CND2X2 U4272 ( .A(n1906), .B(n1905), .Z(n1910) );
  CND2X1 U4273 ( .A(n2085), .B(\m2.addrM64 [1]), .Z(n1912) );
  CND2X1 U4274 ( .A(n2245), .B(\m0.addrM64 [13]), .Z(n2086) );
  CNIVX1 U4275 ( .A(\s1.addr[17] ), .Z(n4095) );
  CNIVX1 U4276 ( .A(\s6.en ), .Z(n4062) );
  CNIVX1 U4277 ( .A(n3378), .Z(n4076) );
  CNIVX1 U4278 ( .A(n4336), .Z(n4094) );
  CNIVX1 U4279 ( .A(\s12.addr[10] ), .Z(n1843) );
  CNIVX1 U4280 ( .A(\s7.addr[16] ), .Z(n4072) );
  CNIVX1 U4281 ( .A(\s8.addr[15] ), .Z(n4109) );
  CNIVX1 U4282 ( .A(n4050), .Z(n4098) );
  CNIVX1 U4283 ( .A(\s1.en ), .Z(n4090) );
  CNIVX1 U4284 ( .A(\s6.en ), .Z(n4075) );
  CNIVX1 U4285 ( .A(\s14.addr[18] ), .Z(n4092) );
  CNIVX1 U4286 ( .A(\s8.en ), .Z(n4085) );
  CNIVX1 U4287 ( .A(\s6.addr [17]), .Z(n1845) );
  CNR2X1 U4288 ( .A(n4258), .B(n3412), .Z(\s13.addr [5]) );
  CNR2X1 U4289 ( .A(n4259), .B(n3405), .Z(\s13.addr [10]) );
  CNR2X1 U4290 ( .A(n3452), .B(n4230), .Z(\s7.addr [22]) );
  CNR2IX1 U4291 ( .B(n5518), .A(n3432), .Z(\m5.ack ) );
  CIVX12 U4292 ( .A(n3445), .Z(\s4.addr [19]) );
  CNR2IX1 U4293 ( .B(n5518), .A(n3439), .Z(\m4.ack ) );
  CAN2X1 U4294 ( .A(n3431), .B(n5518), .Z(\m1.ack ) );
  CAN2X1 U4295 ( .A(n3434), .B(n5518), .Z(\m0.ack ) );
  CNIVX1 U4296 ( .A(n2459), .Z(n3447) );
  CND2X2 U4297 ( .A(n2245), .B(\m0.addrM64 [15]), .Z(n2153) );
  CNR3X2 U4298 ( .A(n2027), .B(n2026), .C(n2025), .Z(n2030) );
  CNIVX1 U4299 ( .A(\c1.sysClk ), .Z(n4386) );
  CND2X2 U4300 ( .A(n2088), .B(\m1.addrM64 [11]), .Z(n1875) );
  CND2X1 U4301 ( .A(n2246), .B(\m6.addrM64 [15]), .Z(n2020) );
  CND2X1 U4302 ( .A(n2088), .B(\m1.addrM64 [15]), .Z(n2157) );
  CIVX2 U4303 ( .A(n2735), .Z(n2140) );
  CNR2IX1 U4304 ( .B(n2165), .A(n2164), .Z(n2169) );
  CNR2X2 U4305 ( .A(n3454), .B(n2171), .Z(n2172) );
  CND2X2 U4306 ( .A(n1993), .B(n1991), .Z(n1895) );
  CND2IX1 U4307 ( .B(n2158), .A(n2157), .Z(n2159) );
  CND2X2 U4308 ( .A(n1994), .B(n1990), .Z(n1896) );
  CND2IX1 U4309 ( .B(n4076), .A(\s10.dbus_out [22]), .Z(n3939) );
  CND2X1 U4310 ( .A(\s2.dbus_out [58]), .B(\s2.addr[16] ), .Z(n1755) );
  CANR2X1 U4311 ( .A(\s7.dbus_out [58]), .B(n4072), .C(\s1.dbus_out [58]), .D(
        n4090), .Z(n1756) );
  CANR2X1 U4312 ( .A(n4099), .B(\s12.dbus_out [58]), .C(\s14.dbus_out [58]), 
        .D(n4092), .Z(n1757) );
  CANR2X1 U4313 ( .A(\s4.dbus_out [58]), .B(n4077), .C(\s5.dbus_out [58]), .D(
        n4078), .Z(n1758) );
  CAOR2X1 U4314 ( .A(\s0.dbus_out [58]), .B(n4083), .C(\s9.addr[16] ), .D(
        \s9.dbus_out [58]), .Z(n1759) );
  CANR1XL U4315 ( .A(\s11.addr[17] ), .B(\s11.dbus_out [58]), .C(n1759), .Z(
        n1760) );
  CANR2X1 U4316 ( .A(data_stm_d[58]), .B(\c1.Breset ), .C(\s6.dbus_out [58]), 
        .D(n4075), .Z(n1761) );
  CANR2X1 U4317 ( .A(\s3.dbus_out [58]), .B(\s3.addr[9] ), .C(
        \s10.dbus_out [58]), .D(n4098), .Z(n1762) );
  CANR2X1 U4318 ( .A(\s8.dbus_out [58]), .B(n4085), .C(\s13.dbus_out [58]), 
        .D(n4110), .Z(n1763) );
  CND8X1 U4319 ( .A(n1755), .B(n1756), .C(n1757), .D(n1758), .E(n1760), .F(
        n1761), .G(n1762), .H(n1763), .Z(n1696) );
  CND2IX1 U4320 ( .B(n4076), .A(\s10.dbus_out [29]), .Z(n4082) );
  CND2X1 U4321 ( .A(\s2.dbus_out [26]), .B(\s2.addr[16] ), .Z(n1764) );
  CANR2X1 U4322 ( .A(\s7.dbus_out [26]), .B(\s7.addr[19] ), .C(
        \s1.dbus_out [26]), .D(n4095), .Z(n1765) );
  CANR2X1 U4323 ( .A(data_stm_d[26]), .B(\c1.Breset ), .C(\s6.dbus_out [26]), 
        .D(n4075), .Z(n1766) );
  CANR2X1 U4324 ( .A(\s8.dbus_out [26]), .B(n4085), .C(\s13.dbus_out [26]), 
        .D(n4110), .Z(n1767) );
  CAN8X1 U4325 ( .A(n1764), .B(n1765), .C(n1766), .D(n3599), .E(n3600), .F(
        n3601), .G(n3602), .H(n1767), .Z(n1768) );
  CANR1XL U4326 ( .A(n4093), .B(\s11.dbus_out [26]), .C(n3603), .Z(n1769) );
  CND2X1 U4327 ( .A(n1768), .B(n1769), .Z(n1728) );
  CND2X1 U4328 ( .A(\s2.dbus_out [59]), .B(\s2.addr[19] ), .Z(n1770) );
  CANR2X1 U4329 ( .A(\s7.dbus_out [59]), .B(n4072), .C(\s1.dbus_out [59]), .D(
        n4090), .Z(n1771) );
  CANR2X1 U4330 ( .A(n4099), .B(\s12.dbus_out [59]), .C(\s14.dbus_out [59]), 
        .D(n4100), .Z(n1772) );
  CANR2X1 U4331 ( .A(\s4.dbus_out [59]), .B(n4077), .C(\s5.dbus_out [59]), .D(
        n4078), .Z(n1773) );
  CAOR2X1 U4332 ( .A(\s0.dbus_out [59]), .B(\s0.en ), .C(\s9.addr[16] ), .D(
        \s9.dbus_out [59]), .Z(n1774) );
  CANR1XL U4333 ( .A(\s11.dbus_out [59]), .B(n4093), .C(n1774), .Z(n1775) );
  CANR2X1 U4334 ( .A(data_stm_d[59]), .B(\c1.Breset ), .C(\s6.dbus_out [59]), 
        .D(n1845), .Z(n1776) );
  CANR2X1 U4335 ( .A(\s3.dbus_out [59]), .B(\s3.addr[9] ), .C(
        \s10.dbus_out [59]), .D(n4098), .Z(n1777) );
  CANR2X1 U4336 ( .A(\s8.dbus_out [59]), .B(n4109), .C(\s13.dbus_out [59]), 
        .D(n4110), .Z(n1778) );
  CND8X1 U4337 ( .A(n1770), .B(n1771), .C(n1772), .D(n1773), .E(n1775), .F(
        n1776), .G(n1777), .H(n1778), .Z(n1695) );
  CIVX1 U4338 ( .A(n2248), .Z(n1779) );
  CANR2X1 U4339 ( .A(n2245), .B(\m0.addrM64 [18]), .C(\m5.addrM64 [18]), .D(
        n1779), .Z(n2051) );
  CND2IX1 U4340 ( .B(n4076), .A(\s10.dbus_out [52]), .Z(n3620) );
  CND2X1 U4341 ( .A(\s2.dbus_out [33]), .B(\s2.addr[19] ), .Z(n1780) );
  CANR2X1 U4342 ( .A(\s7.dbus_out [33]), .B(\s7.addr[19] ), .C(
        \s1.dbus_out [33]), .D(n4090), .Z(n1781) );
  CANR2X1 U4343 ( .A(n4099), .B(\s12.dbus_out [33]), .C(\s14.dbus_out [33]), 
        .D(n4092), .Z(n1782) );
  CANR2X1 U4344 ( .A(\s4.dbus_out [33]), .B(n4091), .C(\s5.dbus_out [33]), .D(
        n4078), .Z(n1783) );
  CAOR2X1 U4345 ( .A(\s0.dbus_out [33]), .B(\s0.addr [13]), .C(\s9.addr [15]), 
        .D(\s9.dbus_out [33]), .Z(n1784) );
  CANR1XL U4346 ( .A(\s11.dbus_out [33]), .B(n4093), .C(n1784), .Z(n1785) );
  CANR2X1 U4347 ( .A(data_stm_d[33]), .B(\c1.Breset ), .C(\s6.dbus_out [33]), 
        .D(\s6.addr [17]), .Z(n1786) );
  CANR2X1 U4348 ( .A(\s3.dbus_out [33]), .B(\s3.addr [18]), .C(
        \s10.dbus_out [33]), .D(\s10.addr[9] ), .Z(n1787) );
  CANR2X1 U4349 ( .A(\s8.dbus_out [33]), .B(\s8.en ), .C(\s13.dbus_out [33]), 
        .D(n4110), .Z(n1788) );
  CND8X1 U4350 ( .A(n1780), .B(n1781), .C(n1782), .D(n1783), .E(n1785), .F(
        n1786), .G(n1787), .H(n1788), .Z(n1721) );
  CND4X1 U4351 ( .A(n2794), .B(n2788), .C(n2789), .D(n2790), .Z(n2797) );
  CANR2X1 U4352 ( .A(n2040), .B(\m3.addrM64 [17]), .C(n2246), .D(
        \m6.addrM64 [17]), .Z(n2044) );
  CIVX1 U4353 ( .A(n3432), .Z(n1789) );
  CAOR2X1 U4354 ( .A(n3435), .B(\m6.DoutM [14]), .C(\m5.DoutM [14]), .D(n1789), 
        .Z(n3150) );
  CIVX2 U4355 ( .A(n3439), .Z(n1790) );
  CAOR2X1 U4356 ( .A(n3436), .B(\m2.DoutM [49]), .C(\m4.DoutM [49]), .D(n1790), 
        .Z(n3026) );
  CANR2X1 U4357 ( .A(n3361), .B(\m3.DoutM [0]), .C(\m1.DoutM [0]), .D(n3431), 
        .Z(n1791) );
  COND3X1 U4358 ( .A(n3432), .B(n2583), .C(n2582), .D(n1791), .Z(n1792) );
  CNR2IXL U4359 ( .B(\m4.DoutM [0]), .A(n3439), .Z(n1793) );
  CNR2X1 U4360 ( .A(n1792), .B(n1793), .Z(n1794) );
  CND3X2 U4361 ( .A(n2580), .B(n2581), .C(n1794), .Z(n4185) );
  CANR2X1 U4362 ( .A(n3361), .B(\m3.DoutM [55]), .C(\m1.DoutM [55]), .D(n3431), 
        .Z(n1795) );
  COND3X1 U4363 ( .A(n3432), .B(n3206), .C(n3205), .D(n1795), .Z(n1796) );
  CNR2IXL U4364 ( .B(\m4.DoutM [55]), .A(n3439), .Z(n1797) );
  CNR2X1 U4365 ( .A(n1796), .B(n1797), .Z(n1798) );
  CND3X2 U4366 ( .A(n3203), .B(n3204), .C(n1798), .Z(n3461) );
  CND2IX1 U4367 ( .B(n4076), .A(\s10.dbus_out [54]), .Z(n3882) );
  CND2X1 U4368 ( .A(\s2.dbus_out [62]), .B(\s2.addr[19] ), .Z(n1799) );
  CANR2X1 U4369 ( .A(\s7.dbus_out [62]), .B(n4336), .C(\s1.dbus_out [62]), .D(
        n4090), .Z(n1800) );
  CANR2X1 U4370 ( .A(n4016), .B(\s12.dbus_out [62]), .C(\s14.dbus_out [62]), 
        .D(\s14.addr [11]), .Z(n1801) );
  CANR2X1 U4371 ( .A(\s4.dbus_out [62]), .B(n4091), .C(\s5.dbus_out [62]), .D(
        n4078), .Z(n1802) );
  CAOR2X1 U4372 ( .A(\s0.dbus_out [62]), .B(n3963), .C(\s9.addr[16] ), .D(
        \s9.dbus_out [62]), .Z(n1803) );
  CANR1XL U4373 ( .A(\s11.dbus_out [62]), .B(n4108), .C(n1803), .Z(n1804) );
  CANR2X1 U4374 ( .A(data_stm_d[62]), .B(\c1.Breset ), .C(\s6.dbus_out [62]), 
        .D(n4075), .Z(n1805) );
  CANR2X1 U4375 ( .A(\s3.dbus_out [62]), .B(\s3.addr[9] ), .C(
        \s10.dbus_out [62]), .D(n4098), .Z(n1806) );
  CANR2X1 U4376 ( .A(\s8.dbus_out [62]), .B(n4085), .C(\s13.dbus_out [62]), 
        .D(n4110), .Z(n1807) );
  CND8X1 U4377 ( .A(n1799), .B(n1800), .C(n1801), .D(n1802), .E(n1804), .F(
        n1805), .G(n1806), .H(n1807), .Z(n1692) );
  CAN3X1 U4378 ( .A(n5518), .B(n1848), .C(n2762), .Z(n2763) );
  CND2IX1 U4379 ( .B(n2078), .A(\m4.addrM64 [17]), .Z(n2042) );
  CNR2IX1 U4380 ( .B(n3409), .A(n2125), .Z(n2781) );
  CAOR2X1 U4381 ( .A(n3431), .B(\m1.DoutM [2]), .C(n3436), .D(\m2.DoutM [2]), 
        .Z(n2444) );
  CIVX1 U4382 ( .A(n3432), .Z(n1808) );
  CAOR2X1 U4383 ( .A(n3435), .B(\m6.DoutM [8]), .C(\m5.DoutM [8]), .D(n1808), 
        .Z(n3032) );
  CIVX1 U4384 ( .A(n3432), .Z(n1809) );
  CAOR2X1 U4385 ( .A(n3231), .B(\m6.DoutM [10]), .C(\m5.DoutM [10]), .D(n1809), 
        .Z(n2269) );
  CIVX1 U4386 ( .A(n3432), .Z(n1810) );
  CAOR2X1 U4387 ( .A(n3435), .B(\m6.DoutM [11]), .C(\m5.DoutM [11]), .D(n1810), 
        .Z(n2652) );
  CAOR2X1 U4388 ( .A(n3434), .B(\m0.DoutM [14]), .C(n3436), .D(\m2.DoutM [14]), 
        .Z(n3151) );
  CAOR2X1 U4389 ( .A(n3431), .B(\m1.DoutM [15]), .C(n3436), .D(\m2.DoutM [15]), 
        .Z(n2993) );
  CIVX1 U4390 ( .A(n3432), .Z(n1811) );
  CAOR2X1 U4391 ( .A(n3435), .B(\m6.DoutM [18]), .C(\m5.DoutM [18]), .D(n1811), 
        .Z(n2260) );
  CAOR2X1 U4392 ( .A(n3435), .B(\m6.DoutM [22]), .C(n3436), .D(\m2.DoutM [22]), 
        .Z(n2702) );
  CAOR2X1 U4393 ( .A(n3431), .B(\m1.DoutM [23]), .C(n3436), .D(\m2.DoutM [23]), 
        .Z(n2328) );
  CIVX1 U4394 ( .A(n3439), .Z(n1812) );
  CAOR2X1 U4395 ( .A(n3436), .B(\m2.DoutM [27]), .C(\m4.DoutM [27]), .D(n1812), 
        .Z(n2872) );
  CIVX1 U4396 ( .A(n3439), .Z(n1813) );
  CAOR2X1 U4397 ( .A(n3436), .B(\m2.DoutM [31]), .C(\m4.DoutM [31]), .D(n1813), 
        .Z(n3080) );
  CIVX1 U4398 ( .A(n3432), .Z(n1814) );
  CAOR2X1 U4399 ( .A(n3435), .B(\m6.DoutM [33]), .C(\m5.DoutM [33]), .D(n1814), 
        .Z(n2356) );
  CAOR2X1 U4400 ( .A(n3431), .B(\m1.DoutM [36]), .C(n3436), .D(\m2.DoutM [36]), 
        .Z(n2987) );
  CAOR2X1 U4401 ( .A(n3434), .B(\m0.DoutM [38]), .C(n3436), .D(\m2.DoutM [38]), 
        .Z(n3235) );
  CAOR2X1 U4402 ( .A(n3431), .B(\m1.DoutM [46]), .C(n3436), .D(\m2.DoutM [46]), 
        .Z(n2414) );
  CIVX1 U4403 ( .A(n3432), .Z(n1815) );
  CAOR2X1 U4404 ( .A(n3435), .B(\m6.DoutM [47]), .C(\m5.DoutM [47]), .D(n1815), 
        .Z(n3368) );
  CIVX1 U4405 ( .A(n3432), .Z(n1816) );
  CAOR2X1 U4406 ( .A(n3435), .B(\m6.DoutM [49]), .C(\m5.DoutM [49]), .D(n1816), 
        .Z(n3027) );
  CIVX1 U4407 ( .A(n3432), .Z(n1817) );
  CAOR2X1 U4408 ( .A(n3435), .B(\m6.DoutM [51]), .C(\m5.DoutM [51]), .D(n1817), 
        .Z(n2473) );
  CIVX1 U4409 ( .A(n3432), .Z(n1818) );
  CAOR2X1 U4410 ( .A(n3435), .B(\m6.DoutM [52]), .C(\m5.DoutM [52]), .D(n1818), 
        .Z(n3313) );
  CAOR2X1 U4411 ( .A(n3435), .B(\m6.DoutM [58]), .C(n3436), .D(\m2.DoutM [58]), 
        .Z(n3199) );
  CAOR2X1 U4412 ( .A(n3434), .B(\m0.DoutM [60]), .C(n3436), .D(\m2.DoutM [60]), 
        .Z(n2686) );
  CIVX1 U4413 ( .A(n3439), .Z(n1819) );
  CAOR2X1 U4414 ( .A(n3436), .B(\m2.DoutM [61]), .C(\m4.DoutM [61]), .D(n1819), 
        .Z(n2679) );
  CIVX1 U4415 ( .A(n3432), .Z(n1820) );
  CAOR2X1 U4416 ( .A(n3435), .B(\m6.addrM64 [20]), .C(\m5.addrM64 [20]), .D(
        n1820), .Z(n2489) );
  CAOR2X1 U4417 ( .A(n3431), .B(\m1.addrM64 [26]), .C(n3436), .D(
        \m2.addrM64 [26]), .Z(n2861) );
  CIVX1 U4418 ( .A(n3432), .Z(n1821) );
  CAOR2X1 U4419 ( .A(n3435), .B(\m6.addrM64 [29]), .C(\m5.addrM64 [29]), .D(
        n1821), .Z(n2321) );
  CAOR2X1 U4420 ( .A(n3435), .B(\m6.addrM64 [32]), .C(n3436), .D(
        \m2.addrM64 [32]), .Z(n3285) );
  CIVX1 U4421 ( .A(n3432), .Z(n1822) );
  CAOR2X1 U4422 ( .A(n3435), .B(\m6.addrM64 [38]), .C(\m5.addrM64 [38]), .D(
        n1822), .Z(n3097) );
  CAOR2X1 U4423 ( .A(n3434), .B(\m0.addrM64 [43]), .C(n3436), .D(
        \m2.addrM64 [43]), .Z(n3010) );
  CIVX1 U4424 ( .A(n3432), .Z(n1823) );
  CAOR2X1 U4425 ( .A(n3435), .B(\m6.addrM64 [45]), .C(\m5.addrM64 [45]), .D(
        n1823), .Z(n3334) );
  CAOR2X1 U4426 ( .A(n3435), .B(\m6.addrM64 [52]), .C(n3436), .D(
        \m2.addrM64 [52]), .Z(n3184) );
  CAOR2X1 U4427 ( .A(n3435), .B(\m6.addrM64 [59]), .C(n3436), .D(
        \m2.addrM64 [59]), .Z(n2943) );
  CAOR2X1 U4428 ( .A(n3435), .B(\m6.addrM64 [63]), .C(n3436), .D(
        \m2.addrM64 [63]), .Z(n3426) );
  CNR2IX1 U4429 ( .B(\m1.addrM64 [2]), .A(n2067), .Z(n2634) );
  CANR2X1 U4430 ( .A(n4090), .B(\s1.dbus_out [9]), .C(n4094), .D(
        \s7.dbus_out [9]), .Z(n1824) );
  CANR2X1 U4431 ( .A(\s6.addr [17]), .B(\s6.dbus_out [9]), .C(data_stm_d[9]), 
        .D(\c1.Breset ), .Z(n1825) );
  CND2X1 U4432 ( .A(n1824), .B(n1825), .Z(n1826) );
  CANR1XL U4433 ( .A(\s2.dbus_out [9]), .B(\s2.addr[19] ), .C(n1826), .Z(n3776) );
  CANR2X1 U4434 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [11]), .C(n4072), .D(
        \s7.dbus_out [11]), .Z(n1827) );
  CANR2X1 U4435 ( .A(\s6.addr [17]), .B(\s6.dbus_out [11]), .C(data_stm_d[11]), 
        .D(\c1.Breset ), .Z(n1828) );
  CND2X1 U4436 ( .A(n1827), .B(n1828), .Z(n1829) );
  CANR1XL U4437 ( .A(\s2.dbus_out [11]), .B(\s2.addr[16] ), .C(n1829), .Z(
        n3756) );
  CND2IX1 U4438 ( .B(n4076), .A(\s10.dbus_out [41]), .Z(n4020) );
  CNR2IX1 U4439 ( .B(n4185), .A(n3251), .Z(\s6.SbusIn [0]) );
  CNR2IX1 U4440 ( .B(n3461), .A(n2812), .Z(\s5.SbusIn [55]) );
  CNR2IX1 U4441 ( .B(n4154), .A(n3453), .Z(\s1.SbusIn [7]) );
  CND2X1 U4442 ( .A(\s2.dbus_out [17]), .B(\s2.addr[16] ), .Z(n1830) );
  CANR2X1 U4443 ( .A(\s7.dbus_out [17]), .B(\s7.en ), .C(\s1.dbus_out [17]), 
        .D(\s1.addr[17] ), .Z(n1831) );
  CANR2X1 U4444 ( .A(n4099), .B(\s12.dbus_out [17]), .C(\s14.dbus_out [17]), 
        .D(n4092), .Z(n1832) );
  CANR2X1 U4445 ( .A(\s4.dbus_out [17]), .B(\s4.addr [19]), .C(
        \s5.dbus_out [17]), .D(n4078), .Z(n1833) );
  CAOR2X1 U4446 ( .A(\s0.dbus_out [17]), .B(\s0.addr [13]), .C(n5590), .D(
        \s9.dbus_out [17]), .Z(n1834) );
  CANR1XL U4447 ( .A(\s11.dbus_out [17]), .B(n4093), .C(n1834), .Z(n1835) );
  CANR2X1 U4448 ( .A(data_stm_d[17]), .B(\c1.Breset ), .C(\s6.dbus_out [17]), 
        .D(n1845), .Z(n1836) );
  CANR2X1 U4449 ( .A(\s3.dbus_out [17]), .B(\s3.addr [18]), .C(
        \s10.dbus_out [17]), .D(\s10.addr[9] ), .Z(n1837) );
  CANR2X1 U4450 ( .A(\s8.dbus_out [17]), .B(n4085), .C(\s13.dbus_out [17]), 
        .D(n4110), .Z(n1838) );
  CND8X1 U4451 ( .A(n1830), .B(n1831), .C(n1832), .D(n1833), .E(n1835), .F(
        n1836), .G(n1837), .H(n1838), .Z(n1737) );
  CIVX8 U4452 ( .A(n2621), .Z(n2456) );
  CND2X2 U4453 ( .A(n2125), .B(n2014), .Z(n2015) );
  CIVX12 U4454 ( .A(n2435), .Z(n3415) );
  CNIVX3 U4455 ( .A(n2223), .Z(n3418) );
  CND2IXL U4456 ( .B(n1911), .A(\m6.addrM64 [1]), .Z(n1914) );
  CND2X2 U4457 ( .A(n2753), .B(n2623), .Z(n1839) );
  CND2X2 U4458 ( .A(n2753), .B(n2623), .Z(n2295) );
  CIVX8 U4459 ( .A(n2045), .Z(n2040) );
  CAN2XL U4460 ( .A(n3413), .B(n4336), .Z(\s7.addr [7]) );
  CAN2XL U4461 ( .A(n4336), .B(n4179), .Z(\s7.addr [33]) );
  CIVX4 U4462 ( .A(n1872), .Z(n2067) );
  CNIVX1 U4463 ( .A(\s12.addr[10] ), .Z(n1840) );
  CND2X1 U4464 ( .A(n2792), .B(n2791), .Z(n2796) );
  CND2X1 U4465 ( .A(n2791), .B(n4257), .Z(n2126) );
  CAN2X2 U4466 ( .A(\m1.addrM64 [18]), .B(n2088), .Z(n1841) );
  CNR2X2 U4467 ( .A(n1841), .B(n2046), .Z(n2053) );
  CIVX20 U4468 ( .A(n3406), .Z(\s14.addr[17] ) );
  CNIVX1 U4469 ( .A(n3090), .Z(n1842) );
  CNIVX4 U4470 ( .A(n2855), .Z(n3090) );
  CIVX16 U4471 ( .A(n3414), .Z(\s12.addr[10] ) );
  CND2X2 U4472 ( .A(n2140), .B(n2755), .Z(n2177) );
  CND2X1 U4473 ( .A(n2108), .B(n2111), .Z(n2006) );
  CAN2X1 U4474 ( .A(\s13.addr[15] ), .B(n4140), .Z(\s13.addr [63]) );
  CND3X1 U4475 ( .A(n3484), .B(n3405), .C(n2288), .Z(n2290) );
  CND3X2 U4476 ( .A(n1952), .B(n1951), .C(n1950), .Z(n1953) );
  CNIVX16 U4477 ( .A(n1968), .Z(n3476) );
  CIVX4 U4478 ( .A(n3476), .Z(n3412) );
  CAN2X1 U4479 ( .A(\m2.addrM64 [14]), .B(n1944), .Z(n2025) );
  CIVX12 U4480 ( .A(n4422), .Z(n1870) );
  CIVX4 U4481 ( .A(n2812), .Z(n1844) );
  CIVX12 U4482 ( .A(n2513), .Z(n4405) );
  CIVX2 U4483 ( .A(n3240), .Z(\s5.addr[14] ) );
  CNIVX1 U4484 ( .A(n2812), .Z(n3240) );
  CNR2X4 U4485 ( .A(n2311), .B(n2310), .Z(n2312) );
  CND2X2 U4486 ( .A(n3384), .B(n3389), .Z(n1858) );
  CND3X1 U4487 ( .A(n2210), .B(n2789), .C(n2209), .Z(n2214) );
  CND3X2 U4488 ( .A(n2791), .B(n2789), .C(n2623), .Z(n2120) );
  CND2X2 U4489 ( .A(n2451), .B(n2450), .Z(n2454) );
  CIVX20 U4490 ( .A(n2455), .Z(\s6.addr [17]) );
  CND3X2 U4491 ( .A(n2789), .B(n2623), .C(n2621), .Z(n2224) );
  CNR2IX1 U4492 ( .B(\m1.addrM64 [0]), .A(n2067), .Z(n1925) );
  CNR2IX1 U4493 ( .B(\m1.addrM64 [14]), .A(n2067), .Z(n2026) );
  CIVX8 U4494 ( .A(n3385), .Z(n1871) );
  CIVX8 U4495 ( .A(n2067), .Z(n2088) );
  CIVDX2 U4496 ( .A(n3385), .Z0(n1859), .Z1(n1846) );
  CIVX3 U4497 ( .A(\m0.ack ), .Z(n3380) );
  CIVDX2 U4498 ( .A(n3409), .Z0(n4257), .Z1(n3456) );
  CIVX3 U4499 ( .A(n3330), .Z(n4110) );
  CIVX2 U4500 ( .A(n1984), .Z(n2167) );
  CIVDX2 U4501 ( .A(n2527), .Z0(n1847), .Z1(n1848) );
  CAN2X1 U4502 ( .A(n4405), .B(n4329), .Z(\s5.SbusIn [6]) );
  CIVX2 U4503 ( .A(n1870), .Z(n3389) );
  CAN2X1 U4504 ( .A(\s9.addr [15]), .B(n4117), .Z(\s9.SbusIn [28]) );
  CAN2X1 U4505 ( .A(\s9.addr [15]), .B(n4151), .Z(\s9.addr [61]) );
  CAN2X1 U4506 ( .A(\s9.addr [15]), .B(n4192), .Z(\s9.SbusIn [2]) );
  CAN2X1 U4507 ( .A(\s9.addr [15]), .B(n3472), .Z(\s9.SbusIn [46]) );
  CND2X4 U4508 ( .A(n1870), .B(n3385), .Z(n1851) );
  CIVX16 U4509 ( .A(n3415), .Z(\s8.addr[15] ) );
  CND2X2 U4510 ( .A(n2782), .B(n2781), .Z(n2800) );
  CND3X1 U4511 ( .A(n2780), .B(n2779), .C(n2778), .Z(n2782) );
  CIVX4 U4512 ( .A(n1870), .Z(n1850) );
  CIVX8 U4513 ( .A(n4419), .Z(n3385) );
  CIVX8 U4514 ( .A(n4420), .Z(n1869) );
  CND3X2 U4515 ( .A(n1850), .B(n3385), .C(n1869), .Z(n1891) );
  CNR2X4 U4516 ( .A(n1851), .B(n1869), .Z(n1944) );
  CANR2X1 U4517 ( .A(n1916), .B(\m5.addrM64 [10]), .C(\m2.addrM64 [10]), .D(
        n1944), .Z(n1853) );
  CIVX8 U4518 ( .A(n1869), .Z(n3384) );
  CNR3X4 U4519 ( .A(n3384), .B(n1870), .C(n3385), .Z(n1882) );
  CNIVX16 U4520 ( .A(n1882), .Z(n2855) );
  CND2X2 U4521 ( .A(n2855), .B(\m3.addrM64 [10]), .Z(n1852) );
  CND2X2 U4522 ( .A(n1853), .B(n1852), .Z(n1856) );
  CND3X2 U4523 ( .A(n1871), .B(n1870), .C(n1869), .Z(n1854) );
  CIVX8 U4524 ( .A(n1854), .Z(n1954) );
  CIVX20 U4525 ( .A(n1954), .Z(n2078) );
  CNR2IX2 U4526 ( .B(\m4.addrM64 [10]), .A(n2078), .Z(n1855) );
  CNR2X4 U4527 ( .A(n1856), .B(n1855), .Z(n1983) );
  CND3X2 U4528 ( .A(n1871), .B(n3384), .C(n1870), .Z(n1857) );
  CIVX8 U4529 ( .A(n1857), .Z(n2057) );
  CND2X1 U4530 ( .A(n2057), .B(\m0.addrM64 [10]), .Z(n1864) );
  CNR2X4 U4531 ( .A(n1858), .B(n1871), .Z(n2247) );
  CND2X1 U4532 ( .A(n2247), .B(\m1.addrM64 [10]), .Z(n1863) );
  CND2X4 U4533 ( .A(n1870), .B(n1869), .Z(n1860) );
  CNR2X4 U4534 ( .A(n1860), .B(n1859), .Z(n1861) );
  CIVX12 U4535 ( .A(n1861), .Z(n1911) );
  CIVX12 U4536 ( .A(n1911), .Z(n1961) );
  CND3X2 U4537 ( .A(n1864), .B(n1863), .C(n1862), .Z(n1865) );
  CIVX4 U4538 ( .A(n1865), .Z(n1982) );
  CND2X4 U4539 ( .A(n1983), .B(n1982), .Z(n2203) );
  CIVX8 U4540 ( .A(n2203), .Z(n2613) );
  CANR2X2 U4541 ( .A(n1961), .B(\m6.addrM64 [11]), .C(\m5.addrM64 [11]), .D(
        n1916), .Z(n1868) );
  CIVX4 U4542 ( .A(n1944), .Z(n1876) );
  CIVX12 U4543 ( .A(n1876), .Z(n2085) );
  CND2X2 U4544 ( .A(n2085), .B(\m2.addrM64 [11]), .Z(n1867) );
  CIVX20 U4545 ( .A(n2078), .Z(n2252) );
  CND2X4 U4546 ( .A(n2252), .B(\m4.addrM64 [11]), .Z(n1866) );
  CND3X4 U4547 ( .A(n1868), .B(n1867), .C(n1866), .Z(n2200) );
  CNR3X4 U4548 ( .A(n1871), .B(n1870), .C(n1869), .Z(n1872) );
  CND2X4 U4549 ( .A(n2855), .B(\m3.addrM64 [11]), .Z(n1874) );
  CND2X1 U4550 ( .A(n2057), .B(\m0.addrM64 [11]), .Z(n1873) );
  CIVX4 U4551 ( .A(n2201), .Z(n2225) );
  CND2X4 U4552 ( .A(n2226), .B(n2225), .Z(n2189) );
  CIVX12 U4553 ( .A(n2057), .Z(n1894) );
  CIVX12 U4554 ( .A(n1894), .Z(n2245) );
  CND2X4 U4555 ( .A(n2245), .B(\m0.addrM64 [8]), .Z(n1881) );
  CNR2IX1 U4556 ( .B(\m2.addrM64 [8]), .A(n1876), .Z(n1877) );
  CIVX2 U4557 ( .A(n1877), .Z(n1880) );
  CNIVX4 U4558 ( .A(n1916), .Z(n2089) );
  CND2X1 U4559 ( .A(n1954), .B(\m4.addrM64 [8]), .Z(n1878) );
  CND4X4 U4560 ( .A(n1881), .B(n1880), .C(n1879), .D(n1878), .Z(n2151) );
  CNIVX4 U4561 ( .A(n1882), .Z(n2018) );
  CNIVX4 U4562 ( .A(n2018), .Z(n2342) );
  CND2X2 U4563 ( .A(n2342), .B(\m3.addrM64 [8]), .Z(n1885) );
  CIVX12 U4564 ( .A(n1911), .Z(n2246) );
  CND3X4 U4565 ( .A(n1885), .B(n1884), .C(n1883), .Z(n2152) );
  CNR2X4 U4566 ( .A(n2151), .B(n2152), .Z(n2199) );
  CNR2IX4 U4567 ( .B(\m4.addrM64 [9]), .A(n2078), .Z(n2164) );
  CIVX2 U4568 ( .A(n2164), .Z(n1886) );
  CNIVX4 U4569 ( .A(n1916), .Z(n2073) );
  CND2X4 U4570 ( .A(n2073), .B(\m5.addrM64 [9]), .Z(n1985) );
  CND2X4 U4571 ( .A(n2855), .B(\m3.addrM64 [9]), .Z(n2165) );
  CND2X4 U4572 ( .A(n2085), .B(\m2.addrM64 [9]), .Z(n1984) );
  CND4X4 U4573 ( .A(n1886), .B(n1985), .C(n2165), .D(n1984), .Z(n2187) );
  CND2X4 U4574 ( .A(n2246), .B(\m6.addrM64 [9]), .Z(n1889) );
  CND2X1 U4575 ( .A(n2247), .B(\m1.addrM64 [9]), .Z(n1888) );
  CND2X1 U4576 ( .A(n2057), .B(\m0.addrM64 [9]), .Z(n1887) );
  CND3X4 U4577 ( .A(n1889), .B(n1888), .C(n1887), .Z(n2188) );
  CNR2X4 U4578 ( .A(n2187), .B(n2188), .Z(n2287) );
  CND4X4 U4579 ( .A(n2613), .B(n2189), .C(n2199), .D(n2287), .Z(n2100) );
  CIVX4 U4580 ( .A(n2100), .Z(n2791) );
  CND2X2 U4581 ( .A(n2088), .B(\m1.addrM64 [3]), .Z(n1997) );
  CND2X4 U4582 ( .A(n2246), .B(\m6.addrM64 [3]), .Z(n1992) );
  CNR2IX2 U4583 ( .B(\m4.addrM64 [3]), .A(n2078), .Z(n1998) );
  CNR2X2 U4584 ( .A(n1890), .B(n1998), .Z(n2144) );
  CIVDX4 U4585 ( .A(n1891), .Z0(n1916), .Z1(n2248) );
  CIVX2 U4586 ( .A(\m5.addrM64 [3]), .Z(n1892) );
  CNR2X4 U4587 ( .A(n2248), .B(n1892), .Z(n1893) );
  CIVX8 U4588 ( .A(n1893), .Z(n1994) );
  CND2X4 U4589 ( .A(n2085), .B(\m2.addrM64 [3]), .Z(n1990) );
  CIVX4 U4590 ( .A(n1894), .Z(n1933) );
  CND2X2 U4591 ( .A(n2855), .B(\m3.addrM64 [3]), .Z(n1991) );
  CNR2X4 U4592 ( .A(n1896), .B(n1895), .Z(n2143) );
  CND2X4 U4593 ( .A(n2144), .B(n2143), .Z(n2099) );
  CND2X2 U4594 ( .A(n2246), .B(\m6.addrM64 [2]), .Z(n1898) );
  CND2X4 U4595 ( .A(n2085), .B(\m2.addrM64 [2]), .Z(n1897) );
  CND2X4 U4596 ( .A(n1898), .B(n1897), .Z(n2635) );
  CNR2X4 U4597 ( .A(n2634), .B(n2635), .Z(n1903) );
  CND2X4 U4598 ( .A(n2245), .B(\m0.addrM64 [2]), .Z(n1900) );
  CND2X4 U4599 ( .A(n2252), .B(\m4.addrM64 [2]), .Z(n1899) );
  CND2X4 U4600 ( .A(n1900), .B(n1899), .Z(n1901) );
  CIVX8 U4601 ( .A(n1901), .Z(n2637) );
  CNIVX1 U4602 ( .A(n1916), .Z(n1904) );
  CNIVX2 U4603 ( .A(n2855), .Z(n1902) );
  CND2X4 U4604 ( .A(n1902), .B(\m3.addrM64 [2]), .Z(n2633) );
  CND4X4 U4605 ( .A(n1903), .B(n2637), .C(n2632), .D(n2633), .Z(n2523) );
  CNR2X4 U4606 ( .A(n2099), .B(n2523), .Z(n2754) );
  CNIVX4 U4607 ( .A(n2018), .Z(n3430) );
  CND2X2 U4608 ( .A(n3430), .B(\m3.addrM64 [1]), .Z(n1906) );
  CND2X1 U4609 ( .A(n1904), .B(\m5.addrM64 [1]), .Z(n1905) );
  CND2X2 U4610 ( .A(n2245), .B(\m0.addrM64 [1]), .Z(n1907) );
  CND2X2 U4611 ( .A(n1908), .B(n1907), .Z(n1909) );
  CNR2X4 U4612 ( .A(n1910), .B(n1909), .Z(n2146) );
  CND2X1 U4613 ( .A(n2247), .B(\m1.addrM64 [1]), .Z(n1913) );
  CAN3X2 U4614 ( .A(n1914), .B(n1913), .C(n1912), .Z(n2145) );
  CND2X4 U4615 ( .A(n2146), .B(n2145), .Z(n2774) );
  CNIVX4 U4616 ( .A(n2855), .Z(n2263) );
  CND2X4 U4617 ( .A(n2263), .B(\m3.addrM64 [0]), .Z(n1915) );
  CIVX4 U4618 ( .A(n1915), .Z(n1921) );
  CND2XL U4619 ( .A(n1916), .B(\m5.addrM64 [0]), .Z(n1919) );
  CND2X1 U4620 ( .A(n2057), .B(\m0.addrM64 [0]), .Z(n1918) );
  CND2X2 U4621 ( .A(n2246), .B(\m6.addrM64 [0]), .Z(n1917) );
  CND3X2 U4622 ( .A(n1919), .B(n1918), .C(n1917), .Z(n1920) );
  CNR2X4 U4623 ( .A(n1921), .B(n1920), .Z(n1927) );
  CND2X4 U4624 ( .A(n2252), .B(\m4.addrM64 [0]), .Z(n1923) );
  CND2X2 U4625 ( .A(n2085), .B(\m2.addrM64 [0]), .Z(n1922) );
  CND2X2 U4626 ( .A(n1923), .B(n1922), .Z(n1924) );
  CNR2X4 U4627 ( .A(n1925), .B(n1924), .Z(n1926) );
  CND2X4 U4628 ( .A(n1927), .B(n1926), .Z(n4337) );
  CND2X2 U4629 ( .A(n2774), .B(n4337), .Z(n1928) );
  CND2X4 U4630 ( .A(n2754), .B(n1928), .Z(n2629) );
  CIVX3 U4631 ( .A(n2629), .Z(n2179) );
  CNIVX4 U4632 ( .A(n1944), .Z(n2244) );
  CND2X2 U4633 ( .A(n2244), .B(\m2.addrM64 [7]), .Z(n1929) );
  CIVX3 U4634 ( .A(n1929), .Z(n1932) );
  CND2X4 U4635 ( .A(n1961), .B(\m6.addrM64 [7]), .Z(n1930) );
  CIVX2 U4636 ( .A(n1930), .Z(n1931) );
  CNR2X4 U4637 ( .A(n1932), .B(n1931), .Z(n1977) );
  CND2X4 U4638 ( .A(n2018), .B(\m3.addrM64 [7]), .Z(n1969) );
  CNR2IX4 U4639 ( .B(\m4.addrM64 [7]), .A(n2078), .Z(n1971) );
  CIVX2 U4640 ( .A(n1971), .Z(n1934) );
  CND2X4 U4641 ( .A(n1933), .B(\m0.addrM64 [7]), .Z(n1973) );
  CNR2IX4 U4642 ( .B(n1969), .A(n1935), .Z(n1938) );
  CND2X4 U4643 ( .A(n2088), .B(\m1.addrM64 [7]), .Z(n1976) );
  CIVX2 U4644 ( .A(n1976), .Z(n1936) );
  CNR2IX4 U4645 ( .B(\m5.addrM64 [7]), .A(n2248), .Z(n1972) );
  CNR2X2 U4646 ( .A(n1936), .B(n1972), .Z(n1937) );
  CND3X4 U4647 ( .A(n1938), .B(n1977), .C(n1937), .Z(n2149) );
  CNR2IX2 U4648 ( .B(\m4.addrM64 [6]), .A(n2078), .Z(n1939) );
  CIVX2 U4649 ( .A(n1939), .Z(n1941) );
  CND2X2 U4650 ( .A(n1961), .B(\m6.addrM64 [6]), .Z(n1940) );
  CND3X4 U4651 ( .A(n1942), .B(n1941), .C(n1940), .Z(n1943) );
  CIVX8 U4652 ( .A(n1943), .Z(n2138) );
  CIVX2 U4653 ( .A(\m5.addrM64 [6]), .Z(n1946) );
  CND2X1 U4654 ( .A(n1944), .B(\m2.addrM64 [6]), .Z(n1945) );
  COND1X2 U4655 ( .A(n1946), .B(n2248), .C(n1945), .Z(n2118) );
  CND2X1 U4656 ( .A(n2057), .B(\m0.addrM64 [6]), .Z(n1947) );
  CND2X2 U4657 ( .A(n1948), .B(n1947), .Z(n2119) );
  CNR2X2 U4658 ( .A(n2118), .B(n2119), .Z(n1949) );
  CND2X4 U4659 ( .A(n2138), .B(n1949), .Z(n2101) );
  CND2X4 U4660 ( .A(n2149), .B(n2101), .Z(n2792) );
  CND2X4 U4661 ( .A(n2088), .B(\m1.addrM64 [5]), .Z(n1952) );
  CND2X4 U4662 ( .A(n2085), .B(\m2.addrM64 [5]), .Z(n1951) );
  CND2X2 U4663 ( .A(n2855), .B(\m3.addrM64 [5]), .Z(n1950) );
  CIVX4 U4664 ( .A(n1953), .Z(n2106) );
  CND2X4 U4665 ( .A(n2073), .B(\m5.addrM64 [5]), .Z(n1957) );
  CND2X1 U4666 ( .A(n1954), .B(\m4.addrM64 [5]), .Z(n1956) );
  CND2X2 U4667 ( .A(n1961), .B(\m6.addrM64 [5]), .Z(n1955) );
  CND3X4 U4668 ( .A(n1957), .B(n1956), .C(n1955), .Z(n2104) );
  CND2X1 U4669 ( .A(n2057), .B(\m0.addrM64 [5]), .Z(n2008) );
  CNR2X4 U4670 ( .A(n2104), .B(n2103), .Z(n1958) );
  CND2X4 U4671 ( .A(n2106), .B(n1958), .Z(n1968) );
  CIVX4 U4672 ( .A(n2018), .Z(n2045) );
  CND2X4 U4673 ( .A(n2040), .B(\m3.addrM64 [4]), .Z(n2003) );
  CND2X2 U4674 ( .A(n2111), .B(n2002), .Z(n1960) );
  CNR2X2 U4675 ( .A(n1960), .B(n1959), .Z(n1965) );
  CND2X4 U4676 ( .A(n2085), .B(\m2.addrM64 [4]), .Z(n1963) );
  CND2X2 U4677 ( .A(n1961), .B(\m6.addrM64 [4]), .Z(n1962) );
  CND2X4 U4678 ( .A(n1963), .B(n1962), .Z(n2004) );
  CIVX2 U4679 ( .A(n2004), .Z(n1964) );
  CND2X4 U4680 ( .A(n2245), .B(\m0.addrM64 [4]), .Z(n2109) );
  CND4X2 U4681 ( .A(n2003), .B(n1965), .C(n1964), .D(n2109), .Z(n1966) );
  CND2X4 U4682 ( .A(n1968), .B(n1966), .Z(n2780) );
  CND2X4 U4683 ( .A(n2792), .B(n2780), .Z(n1980) );
  CIVX2 U4684 ( .A(n1980), .Z(n1967) );
  CND3X2 U4685 ( .A(n2791), .B(n2179), .C(n1967), .Z(n2017) );
  CIVX2 U4686 ( .A(n1969), .Z(n1970) );
  CNR2X2 U4687 ( .A(n1971), .B(n1970), .Z(n1975) );
  CIVX2 U4688 ( .A(n1972), .Z(n1974) );
  CND3X4 U4689 ( .A(n1975), .B(n1974), .C(n1973), .Z(n2117) );
  CND2X4 U4690 ( .A(n1979), .B(n1978), .Z(n3409) );
  CND2X2 U4691 ( .A(n2791), .B(n1981), .Z(n2016) );
  CND2X4 U4692 ( .A(n1983), .B(n1982), .Z(n2208) );
  COND1X2 U4693 ( .A(n2151), .B(n2152), .C(n2208), .Z(n2122) );
  CIVX2 U4694 ( .A(n2189), .Z(n1989) );
  CIVX2 U4695 ( .A(n2188), .Z(n1988) );
  CIVX4 U4696 ( .A(n1985), .Z(n2166) );
  CIVX2 U4697 ( .A(n2165), .Z(n1986) );
  CNR3X2 U4698 ( .A(n2166), .B(n1986), .C(n2164), .Z(n1987) );
  CND2X4 U4699 ( .A(n1989), .B(n2198), .Z(n2123) );
  CNR2X4 U4700 ( .A(n2122), .B(n2123), .Z(n2125) );
  CND4X2 U4701 ( .A(n1993), .B(n1992), .C(n1991), .D(n1990), .Z(n1996) );
  CIVX2 U4702 ( .A(n1994), .Z(n1995) );
  CNR2X2 U4703 ( .A(n1996), .B(n1995), .Z(n2001) );
  CIVX2 U4704 ( .A(n1997), .Z(n1999) );
  CIVX8 U4705 ( .A(n2772), .Z(n3459) );
  CND2X4 U4706 ( .A(n2003), .B(n2002), .Z(n2005) );
  CNR2X4 U4707 ( .A(n2005), .B(n2004), .Z(n2112) );
  CIVX4 U4708 ( .A(n2112), .Z(n2007) );
  CNR2X4 U4709 ( .A(n2007), .B(n2006), .Z(n2543) );
  CIVDX2 U4710 ( .A(n2008), .Z0(n2103), .Z1(n2009) );
  CND2X2 U4711 ( .A(n2109), .B(n2009), .Z(n2010) );
  CIVX2 U4712 ( .A(n2010), .Z(n2011) );
  CND2X2 U4713 ( .A(n2011), .B(n2106), .Z(n2013) );
  CNIVX3 U4714 ( .A(n2104), .Z(n2012) );
  CNR2X4 U4715 ( .A(n2013), .B(n2012), .Z(n2541) );
  CND2X4 U4716 ( .A(n2543), .B(n2541), .Z(n2620) );
  CIVX8 U4717 ( .A(n2620), .Z(n2623) );
  CANR1X2 U4718 ( .A(n3459), .B(n2623), .C(n2792), .Z(n2014) );
  CND3X2 U4719 ( .A(n2017), .B(n2016), .C(n2015), .Z(n2096) );
  CNIVX4 U4720 ( .A(n2018), .Z(n2019) );
  CND2X2 U4721 ( .A(n2019), .B(\m3.addrM64 [15]), .Z(n2021) );
  CND2X4 U4722 ( .A(n2021), .B(n2020), .Z(n2156) );
  CIVX2 U4723 ( .A(n2157), .Z(n2022) );
  CNR2X4 U4724 ( .A(n2156), .B(n2022), .Z(n2131) );
  CND2X2 U4725 ( .A(n2252), .B(\m4.addrM64 [15]), .Z(n2024) );
  CND2X1 U4726 ( .A(n2244), .B(\m2.addrM64 [15]), .Z(n2023) );
  CND2X2 U4727 ( .A(n2024), .B(n2023), .Z(n2158) );
  CAN2X2 U4728 ( .A(n2073), .B(\m5.addrM64 [15]), .Z(n2155) );
  CNR2X4 U4729 ( .A(n2158), .B(n2155), .Z(n2130) );
  CND3X4 U4730 ( .A(n2131), .B(n2153), .C(n2130), .Z(n2761) );
  CNR2IX2 U4731 ( .B(\m4.addrM64 [14]), .A(n2078), .Z(n2027) );
  CANR2X2 U4732 ( .A(n2245), .B(\m0.addrM64 [14]), .C(\m5.addrM64 [14]), .D(
        n2089), .Z(n2029) );
  CANR2X4 U4733 ( .A(n3090), .B(\m3.addrM64 [14]), .C(\m6.addrM64 [14]), .D(
        n2246), .Z(n2028) );
  CND3X4 U4734 ( .A(n2030), .B(n2029), .C(n2028), .Z(n2527) );
  CND2X1 U4735 ( .A(n1847), .B(n5518), .Z(n2031) );
  CNIVX4 U4736 ( .A(n2855), .Z(n3299) );
  CANR2X4 U4737 ( .A(n3299), .B(\m3.addrM64 [19]), .C(\m1.addrM64 [19]), .D(
        n2088), .Z(n2039) );
  CAN2X1 U4738 ( .A(n2252), .B(\m4.addrM64 [19]), .Z(n2035) );
  CND2X2 U4739 ( .A(n2085), .B(\m2.addrM64 [19]), .Z(n2033) );
  CND2X2 U4740 ( .A(n2246), .B(\m6.addrM64 [19]), .Z(n2032) );
  CND2X2 U4741 ( .A(n2033), .B(n2032), .Z(n2034) );
  CNR2X2 U4742 ( .A(n2035), .B(n2034), .Z(n2038) );
  CANR1X2 U4743 ( .A(n2245), .B(\m0.addrM64 [19]), .C(n2036), .Z(n2037) );
  CND3X4 U4744 ( .A(n2039), .B(n2038), .C(n2037), .Z(n2056) );
  CANR2X1 U4745 ( .A(n2088), .B(\m1.addrM64 [17]), .C(\m2.addrM64 [17]), .D(
        n2085), .Z(n2043) );
  CND4X2 U4746 ( .A(n2044), .B(n2043), .C(n2042), .D(n2041), .Z(n2055) );
  CNR2IX2 U4747 ( .B(\m3.addrM64 [18]), .A(n2045), .Z(n2046) );
  CND2X1 U4748 ( .A(n2244), .B(\m2.addrM64 [18]), .Z(n2047) );
  CND3X2 U4749 ( .A(n2053), .B(n2052), .C(n2051), .Z(n2054) );
  CND3X4 U4750 ( .A(n2056), .B(n2054), .C(n2055), .Z(n2233) );
  CIVX8 U4751 ( .A(n2233), .Z(n2465) );
  CND2X1 U4752 ( .A(n2057), .B(\m0.addrM64 [16]), .Z(n2061) );
  CIVX2 U4753 ( .A(\m6.addrM64 [16]), .Z(n2058) );
  CNR2X4 U4754 ( .A(n2059), .B(n2058), .Z(n2060) );
  CNR2IX2 U4755 ( .B(n2061), .A(n2060), .Z(n2065) );
  CNR2IX2 U4756 ( .B(\m5.addrM64 [16]), .A(n2248), .Z(n2063) );
  CNR2IX2 U4757 ( .B(\m4.addrM64 [16]), .A(n2078), .Z(n2062) );
  CNR2X4 U4758 ( .A(n2063), .B(n2062), .Z(n2064) );
  CND2X2 U4759 ( .A(n2065), .B(n2064), .Z(n2066) );
  CIVX3 U4760 ( .A(n2066), .Z(n2070) );
  CANR2X2 U4761 ( .A(n3299), .B(\m3.addrM64 [16]), .C(\m2.addrM64 [16]), .D(
        n2085), .Z(n2069) );
  CND3X4 U4762 ( .A(n2070), .B(n2069), .C(n2068), .Z(n2552) );
  CIVX2 U4763 ( .A(n2245), .Z(n2072) );
  CIVX2 U4764 ( .A(\m0.addrM64 [12]), .Z(n2071) );
  CNR2X2 U4765 ( .A(n2072), .B(n2071), .Z(n2077) );
  CND2X2 U4766 ( .A(n2073), .B(\m5.addrM64 [12]), .Z(n2074) );
  CND2X2 U4767 ( .A(n2075), .B(n2074), .Z(n2076) );
  CNR2X4 U4768 ( .A(n2077), .B(n2076), .Z(n2184) );
  CNR2IX2 U4769 ( .B(\m4.addrM64 [12]), .A(n2078), .Z(n2079) );
  CIVX2 U4770 ( .A(n2079), .Z(n2080) );
  CND2X2 U4771 ( .A(n2081), .B(n2080), .Z(n2185) );
  CIVX2 U4772 ( .A(n2185), .Z(n2082) );
  CNIVX4 U4773 ( .A(n2855), .Z(n3137) );
  CND2X4 U4774 ( .A(n3137), .B(\m3.addrM64 [12]), .Z(n2183) );
  CND3X2 U4775 ( .A(n2184), .B(n2082), .C(n2183), .Z(n2083) );
  CND2X4 U4776 ( .A(n2552), .B(n2083), .Z(n2084) );
  CIVX8 U4777 ( .A(n2084), .Z(n2783) );
  CANR2X2 U4778 ( .A(n2252), .B(\m4.addrM64 [13]), .C(\m2.addrM64 [13]), .D(
        n2085), .Z(n2087) );
  CND2X2 U4779 ( .A(n2087), .B(n2086), .Z(n2163) );
  CANR2X4 U4780 ( .A(n2088), .B(\m1.addrM64 [13]), .C(\m6.addrM64 [13]), .D(
        n2246), .Z(n2092) );
  CND2X2 U4781 ( .A(n2089), .B(\m5.addrM64 [13]), .Z(n2091) );
  CND2X1 U4782 ( .A(n2855), .B(\m3.addrM64 [13]), .Z(n2090) );
  CND3X4 U4783 ( .A(n2092), .B(n2091), .C(n2090), .Z(n2162) );
  CNR2X2 U4784 ( .A(n2163), .B(n2162), .Z(n2232) );
  CIVX2 U4785 ( .A(n2232), .Z(n2093) );
  CNR2X2 U4786 ( .A(n2094), .B(n2129), .Z(n2095) );
  CND2X4 U4787 ( .A(n2096), .B(n2095), .Z(n2097) );
  CIVX8 U4788 ( .A(n2097), .Z(n2098) );
  CIVX16 U4789 ( .A(n2098), .Z(n3451) );
  CIVX8 U4790 ( .A(n3451), .Z(\s7.addr[16] ) );
  CIVX8 U4791 ( .A(n3451), .Z(\s7.addr[19] ) );
  CND2X4 U4792 ( .A(n2523), .B(n2099), .Z(n2621) );
  CNR2X2 U4793 ( .A(n2100), .B(n2456), .Z(n2115) );
  CNR2X2 U4794 ( .A(n2116), .B(n2117), .Z(n2102) );
  CNR2X4 U4795 ( .A(n2102), .B(n2101), .Z(n2113) );
  CNR2X2 U4796 ( .A(n2104), .B(n2103), .Z(n2105) );
  CND2X1 U4797 ( .A(n2106), .B(n2105), .Z(n2107) );
  CIVX2 U4798 ( .A(n2107), .Z(n2141) );
  CND4X4 U4799 ( .A(n2112), .B(n2111), .C(n2110), .D(n2109), .Z(n4338) );
  CND3X2 U4800 ( .A(n2113), .B(n2141), .C(n4338), .Z(n2114) );
  CIVX4 U4801 ( .A(n2114), .Z(n2547) );
  CND3X2 U4802 ( .A(n2774), .B(n4337), .C(n2772), .Z(n2230) );
  CND3X2 U4803 ( .A(n2115), .B(n2547), .C(n2230), .Z(n2121) );
  CNR2X4 U4804 ( .A(n2117), .B(n2116), .Z(n2142) );
  CNR2X4 U4805 ( .A(n2119), .B(n2118), .Z(n2137) );
  CND2X4 U4806 ( .A(n2137), .B(n2138), .Z(n2631) );
  CNR2X4 U4807 ( .A(n2142), .B(n2631), .Z(n2789) );
  CND2X4 U4808 ( .A(n2121), .B(n2120), .Z(n2314) );
  CIVX4 U4809 ( .A(n2314), .Z(n2135) );
  CNR2X4 U4810 ( .A(n2123), .B(n2122), .Z(n2794) );
  CIVX4 U4811 ( .A(n2754), .Z(n2790) );
  CND3X4 U4812 ( .A(n2794), .B(n2790), .C(n3476), .Z(n2311) );
  CIVX4 U4813 ( .A(n2792), .Z(n2793) );
  CNR2X4 U4814 ( .A(n2774), .B(n4337), .Z(n2124) );
  CND2X4 U4815 ( .A(n2124), .B(n3459), .Z(n2639) );
  CND2X2 U4816 ( .A(n2793), .B(n2639), .Z(n2310) );
  CNR2X2 U4817 ( .A(n2311), .B(n2310), .Z(n2128) );
  CND2X2 U4818 ( .A(n2127), .B(n2126), .Z(n2313) );
  CNR2X2 U4819 ( .A(n2128), .B(n2313), .Z(n2134) );
  CIVX2 U4820 ( .A(n2129), .Z(n2133) );
  CIVX2 U4821 ( .A(n1848), .Z(n2728) );
  CND3X2 U4822 ( .A(n2131), .B(n2153), .C(n2130), .Z(n2729) );
  CND2X1 U4823 ( .A(n2729), .B(n5518), .Z(n2785) );
  CNR2X2 U4824 ( .A(n2728), .B(n2785), .Z(n2132) );
  CND2X4 U4825 ( .A(n2133), .B(n2132), .Z(n2315) );
  CANR1X4 U4826 ( .A(n2135), .B(n2134), .C(n2315), .Z(n2136) );
  CIVX8 U4827 ( .A(n2136), .Z(n3038) );
  CIVX16 U4828 ( .A(n3038), .Z(\s11.addr[17] ) );
  CIVX8 U4829 ( .A(n2149), .Z(n2542) );
  CND2X2 U4830 ( .A(n2138), .B(n2137), .Z(n2470) );
  CND2X4 U4831 ( .A(n2542), .B(n2139), .Z(n2291) );
  CIVX8 U4832 ( .A(n2291), .Z(n2753) );
  CIVX8 U4833 ( .A(n2753), .Z(n2538) );
  CND2X4 U4834 ( .A(n2538), .B(n4335), .Z(n2735) );
  CND2X2 U4835 ( .A(n2623), .B(n2542), .Z(n2755) );
  CAN2X2 U4836 ( .A(n2142), .B(n2141), .Z(n2736) );
  CND2X2 U4837 ( .A(n2144), .B(n2143), .Z(n2773) );
  CNR2X2 U4838 ( .A(n4337), .B(n2773), .Z(n2750) );
  CND2X2 U4839 ( .A(n2146), .B(n2145), .Z(n3047) );
  CND3X1 U4840 ( .A(n2736), .B(n2750), .C(n3468), .Z(n2147) );
  CNR2X2 U4841 ( .A(n2629), .B(n2147), .Z(n2176) );
  CNR2X2 U4842 ( .A(n3468), .B(n2621), .Z(n2148) );
  CND2X2 U4843 ( .A(n2148), .B(n2547), .Z(n2727) );
  CNIVX4 U4844 ( .A(n2149), .Z(n3413) );
  CND2X4 U4845 ( .A(n3413), .B(n3476), .Z(n2150) );
  CND2X4 U4846 ( .A(n2150), .B(n2792), .Z(n2537) );
  CIVX2 U4847 ( .A(n2537), .Z(n2724) );
  CNR2X4 U4848 ( .A(n2152), .B(n2151), .Z(n2459) );
  CND3X4 U4849 ( .A(n2727), .B(n2724), .C(n3447), .Z(n2175) );
  CND2X4 U4850 ( .A(n2465), .B(n2783), .Z(n2732) );
  CIVX2 U4851 ( .A(n2153), .Z(n2154) );
  CNR3X2 U4852 ( .A(n2156), .B(n2155), .C(n2154), .Z(n2161) );
  CNR2X2 U4853 ( .A(n2159), .B(\c1.Breset ), .Z(n2160) );
  CND3X4 U4854 ( .A(n2527), .B(n2161), .C(n2160), .Z(n2235) );
  CNR2X4 U4855 ( .A(n2163), .B(n2162), .Z(n2731) );
  CNR2X2 U4856 ( .A(n2167), .B(n2166), .Z(n2168) );
  CND2X2 U4857 ( .A(n2169), .B(n2168), .Z(n2170) );
  CNR2X4 U4858 ( .A(n2170), .B(n2188), .Z(n3454) );
  CNR2X1 U4859 ( .A(n2201), .B(n2200), .Z(n2171) );
  CND3X2 U4860 ( .A(n2731), .B(n2172), .C(n2208), .Z(n2173) );
  CNR3X4 U4861 ( .A(n2732), .B(n2235), .C(n2173), .Z(n2174) );
  COND3X4 U4862 ( .A(n2177), .B(n2176), .C(n2175), .D(n2174), .Z(n3407) );
  CIVX4 U4863 ( .A(n3407), .Z(\s12.addr [19]) );
  CIVX8 U4864 ( .A(\s12.addr [19]), .Z(n3414) );
  CIVX12 U4865 ( .A(n3451), .Z(\s7.en ) );
  CAN2X1 U4866 ( .A(n2736), .B(n3478), .Z(n2178) );
  CND2X2 U4867 ( .A(n2179), .B(n2178), .Z(n2450) );
  CAN2X1 U4868 ( .A(n2542), .B(n2631), .Z(n2180) );
  CIVX2 U4869 ( .A(n3476), .Z(n4253) );
  CNR2X1 U4870 ( .A(n4253), .B(n2291), .Z(n2181) );
  CNR2IX2 U4871 ( .B(n2182), .A(n2181), .Z(n2451) );
  CND2X2 U4872 ( .A(n2184), .B(n2183), .Z(n2186) );
  CNR2X4 U4873 ( .A(n2186), .B(n2185), .Z(n2462) );
  CIVX3 U4874 ( .A(n2731), .Z(n2784) );
  CND3X4 U4875 ( .A(n2462), .B(n1847), .C(n2784), .Z(n2614) );
  CIVX2 U4876 ( .A(n2614), .Z(n2191) );
  CND2X2 U4877 ( .A(n2190), .B(n2189), .Z(n2211) );
  CNR2X2 U4878 ( .A(n2211), .B(n2459), .Z(n2618) );
  CND2X2 U4879 ( .A(n2191), .B(n2618), .Z(n2192) );
  CIVX2 U4880 ( .A(n2192), .Z(n2196) );
  CAN2X1 U4881 ( .A(n2208), .B(n5518), .Z(n2193) );
  CND3X1 U4882 ( .A(n2464), .B(n2729), .C(n2193), .Z(n2194) );
  CIVX8 U4883 ( .A(n2465), .Z(n2786) );
  CNR2X2 U4884 ( .A(n2194), .B(n2786), .Z(n2195) );
  CANR1X4 U4885 ( .A(n2450), .B(n2451), .C(n2452), .Z(n2197) );
  CIVX8 U4886 ( .A(n2197), .Z(n3251) );
  CIVX20 U4887 ( .A(n3251), .Z(\s6.en ) );
  CND3X2 U4888 ( .A(n2639), .B(n2790), .C(n4334), .Z(n2207) );
  CND2X4 U4889 ( .A(n2199), .B(n2198), .Z(n2529) );
  CNR2X2 U4890 ( .A(n2291), .B(n2529), .Z(n2206) );
  CIVDX3 U4891 ( .A(n2200), .Z0(n2226), .Z1(n2202) );
  CNR2X2 U4892 ( .A(n2202), .B(n2201), .Z(n3448) );
  CIVX4 U4893 ( .A(n2203), .Z(n3405) );
  CND3X2 U4894 ( .A(n3412), .B(n3484), .C(n3405), .Z(n2204) );
  CIVX2 U4895 ( .A(n2204), .Z(n2205) );
  CND3X2 U4896 ( .A(n2207), .B(n2206), .C(n2205), .Z(n2215) );
  CNR2X1 U4897 ( .A(n2211), .B(n2621), .Z(n2210) );
  CNR3X2 U4898 ( .A(n2459), .B(n2780), .C(n2208), .Z(n2209) );
  CIVX2 U4899 ( .A(n2211), .Z(n2212) );
  CND4X2 U4900 ( .A(n2793), .B(n3405), .C(n2212), .D(n4335), .Z(n2213) );
  CND3X2 U4901 ( .A(n2215), .B(n2214), .C(n2213), .Z(n2221) );
  CND3X2 U4902 ( .A(n2527), .B(n2731), .C(n2761), .Z(n2216) );
  CIVX2 U4903 ( .A(n2216), .Z(n2217) );
  CNR2X4 U4904 ( .A(n2218), .B(n2786), .Z(n2647) );
  CND2X2 U4905 ( .A(n2647), .B(n5518), .Z(n2219) );
  CIVX3 U4906 ( .A(n2219), .Z(n2220) );
  CND2X4 U4907 ( .A(n2221), .B(n2220), .Z(n2222) );
  CIVX12 U4908 ( .A(n2222), .Z(n2435) );
  CIVX8 U4909 ( .A(n2435), .Z(n2223) );
  CND2X2 U4910 ( .A(n2224), .B(n3409), .Z(n2241) );
  CND2X2 U4911 ( .A(n2226), .B(n2225), .Z(n2240) );
  CNR2X4 U4912 ( .A(n2240), .B(n2287), .Z(n2228) );
  CIVX3 U4913 ( .A(n2459), .Z(n2227) );
  CND3X4 U4914 ( .A(n2228), .B(n2227), .C(n2613), .Z(n2645) );
  CIVX2 U4915 ( .A(n2645), .Z(n2229) );
  COND1X2 U4916 ( .A(n4257), .B(n2230), .C(n2229), .Z(n2231) );
  CND2X2 U4917 ( .A(n2241), .B(n2231), .Z(n2239) );
  CND2X2 U4918 ( .A(n2462), .B(n2232), .Z(n2234) );
  CNR2X2 U4919 ( .A(n2234), .B(n2233), .Z(n2237) );
  CIVX3 U4920 ( .A(n2235), .Z(n2467) );
  CIVDX1 U4921 ( .A(n2552), .Z0(n2464), .Z1(n2236) );
  CND3X4 U4922 ( .A(n2237), .B(n2467), .C(n2236), .Z(n2238) );
  CIVX4 U4923 ( .A(n2238), .Z(n2286) );
  CND2X4 U4924 ( .A(n2239), .B(n2286), .Z(n2744) );
  CIVX4 U4925 ( .A(n2240), .Z(n2762) );
  CND2X4 U4926 ( .A(n2613), .B(n2762), .Z(n2528) );
  CNR2X4 U4927 ( .A(n2528), .B(n2529), .Z(n2548) );
  CNR2X2 U4928 ( .A(n2241), .B(n2548), .Z(n2743) );
  CNR2X4 U4929 ( .A(n2744), .B(n2743), .Z(n2242) );
  CIVX8 U4930 ( .A(n2242), .Z(n2243) );
  CIVX20 U4931 ( .A(n2243), .Z(\s3.addr[14] ) );
  CNIVX12 U4932 ( .A(n2244), .Z(n3436) );
  CAN2X1 U4933 ( .A(n3436), .B(n5518), .Z(\m2.ack ) );
  CNIVX12 U4934 ( .A(n2245), .Z(n3434) );
  CIVDX2 U4935 ( .A(n2246), .Z0(n2059), .Z1(n3231) );
  CNIVX20 U4936 ( .A(n3231), .Z(n3435) );
  CAN2X1 U4937 ( .A(n3435), .B(n5518), .Z(\m6.ack ) );
  CIVX16 U4938 ( .A(n3414), .Z(\s12.addr[11] ) );
  CANR2X1 U4939 ( .A(n3431), .B(\m1.DoutM [48]), .C(\m3.DoutM [48]), .D(n3430), 
        .Z(n2257) );
  CNIVX12 U4940 ( .A(n2248), .Z(n3432) );
  CNR2IX1 U4941 ( .B(\m5.DoutM [48]), .A(n3432), .Z(n2249) );
  CANR1X1 U4942 ( .A(n3434), .B(\m0.DoutM [48]), .C(n2249), .Z(n2256) );
  CND2XL U4943 ( .A(n3435), .B(\m6.DoutM [48]), .Z(n2251) );
  CND2XL U4944 ( .A(n3436), .B(\m2.DoutM [48]), .Z(n2250) );
  CND2X1 U4945 ( .A(n2251), .B(n2250), .Z(n2254) );
  CNIVX4 U4946 ( .A(n2252), .Z(n3424) );
  CIVX8 U4947 ( .A(n3424), .Z(n3439) );
  CNR2IX1 U4948 ( .B(\m4.DoutM [48]), .A(n3439), .Z(n2253) );
  CNR2X2 U4949 ( .A(n2254), .B(n2253), .Z(n2255) );
  CND3X4 U4950 ( .A(n2257), .B(n2256), .C(n2255), .Z(n4121) );
  CAN2X1 U4951 ( .A(\s12.addr[11] ), .B(n4121), .Z(\s12.SbusIn [48]) );
  CND2X1 U4952 ( .A(n3434), .B(\m0.DoutM [18]), .Z(n2259) );
  CND2X1 U4953 ( .A(n3436), .B(\m2.DoutM [18]), .Z(n2258) );
  CND2X1 U4954 ( .A(n2259), .B(n2258), .Z(n2261) );
  CNR2X1 U4955 ( .A(n2261), .B(n2260), .Z(n2266) );
  CNR2IX1 U4956 ( .B(\m4.DoutM [18]), .A(n3439), .Z(n2262) );
  CANR1X1 U4957 ( .A(n3431), .B(\m1.DoutM [18]), .C(n2262), .Z(n2265) );
  CNIVX1 U4958 ( .A(n2263), .Z(n3371) );
  CND2X2 U4959 ( .A(n3371), .B(\m3.DoutM [18]), .Z(n2264) );
  CND3X2 U4960 ( .A(n2266), .B(n2265), .C(n2264), .Z(n4180) );
  CAN2XL U4961 ( .A(\s12.addr[11] ), .B(n4180), .Z(\s12.SbusIn [18]) );
  CND2X1 U4962 ( .A(n3434), .B(\m0.DoutM [10]), .Z(n2268) );
  CND2XL U4963 ( .A(n3436), .B(\m2.DoutM [10]), .Z(n2267) );
  CND2X1 U4964 ( .A(n2268), .B(n2267), .Z(n2270) );
  CNR2X1 U4965 ( .A(n2270), .B(n2269), .Z(n2274) );
  CNR2IX1 U4966 ( .B(\m4.DoutM [10]), .A(n3439), .Z(n2271) );
  CANR1X1 U4967 ( .A(n3431), .B(\m1.DoutM [10]), .C(n2271), .Z(n2273) );
  CNIVX2 U4968 ( .A(n3090), .Z(n3361) );
  CND2X1 U4969 ( .A(n3361), .B(\m3.DoutM [10]), .Z(n2272) );
  CND3X2 U4970 ( .A(n2274), .B(n2273), .C(n2272), .Z(n4115) );
  CAN2XL U4971 ( .A(\s12.addr[11] ), .B(n4115), .Z(\s12.SbusIn [10]) );
  CND2XL U4972 ( .A(n3431), .B(\m1.DoutM [3]), .Z(n2276) );
  CND2XL U4973 ( .A(n3436), .B(\m2.DoutM [3]), .Z(n2275) );
  CND2X1 U4974 ( .A(n2276), .B(n2275), .Z(n2278) );
  CNR2IX1 U4975 ( .B(\m4.DoutM [3]), .A(n3439), .Z(n2277) );
  CNR2X1 U4976 ( .A(n2278), .B(n2277), .Z(n2282) );
  CNIVX4 U4977 ( .A(n3137), .Z(n3420) );
  CANR2X1 U4978 ( .A(n3435), .B(\m6.DoutM [3]), .C(\m3.DoutM [3]), .D(n3420), 
        .Z(n2281) );
  CNR2IX1 U4979 ( .B(\m5.DoutM [3]), .A(n3432), .Z(n2279) );
  CAN2XL U4980 ( .A(\s12.addr[10] ), .B(n4200), .Z(\s12.SbusIn [3]) );
  CIVX2 U4981 ( .A(n2529), .Z(n2765) );
  CIVX2 U4982 ( .A(n3405), .Z(n3475) );
  CNR2X2 U4983 ( .A(n3475), .B(n3448), .Z(n2283) );
  CND2X1 U4984 ( .A(n2765), .B(n2283), .Z(n2284) );
  CND2X2 U4985 ( .A(n1839), .B(n2284), .Z(n2285) );
  CND2X4 U4986 ( .A(n2286), .B(n2285), .Z(n2298) );
  CNR2X1 U4987 ( .A(n2459), .B(n2287), .Z(n2288) );
  CNR2X1 U4988 ( .A(n3468), .B(n2621), .Z(n2289) );
  CNR2X2 U4989 ( .A(n2290), .B(n2289), .Z(n2296) );
  CND2X2 U4990 ( .A(n4337), .B(n2773), .Z(n2775) );
  CNR2IX2 U4991 ( .B(n2775), .A(n2291), .Z(n2293) );
  CNR2X2 U4992 ( .A(n2456), .B(n3476), .Z(n2292) );
  CND2X1 U4993 ( .A(n2773), .B(n2774), .Z(n2622) );
  CND4X4 U4994 ( .A(n2295), .B(n2293), .C(n2292), .D(n2622), .Z(n2294) );
  COND1X4 U4995 ( .A(n2296), .B(n1839), .C(n2294), .Z(n2299) );
  CNR2X4 U4996 ( .A(n2298), .B(n2299), .Z(n2297) );
  CIVX8 U4997 ( .A(n2297), .Z(n3406) );
  CNR2X4 U4998 ( .A(n2299), .B(n2298), .Z(n2300) );
  CIVX8 U4999 ( .A(n2300), .Z(n2301) );
  CIVX16 U5000 ( .A(n2301), .Z(\s14.addr[18] ) );
  CND2X1 U5001 ( .A(n3431), .B(\m1.addrM64 [61]), .Z(n2303) );
  CND2XL U5002 ( .A(n3436), .B(\m2.addrM64 [61]), .Z(n2302) );
  CND2X1 U5003 ( .A(n2303), .B(n2302), .Z(n2305) );
  CAN2XL U5004 ( .A(n3424), .B(\m4.addrM64 [61]), .Z(n2304) );
  CNR2X1 U5005 ( .A(n2305), .B(n2304), .Z(n2309) );
  CANR2X1 U5006 ( .A(n3371), .B(\m3.addrM64 [61]), .C(\m6.addrM64 [61]), .D(
        n3435), .Z(n2308) );
  CNR2IX1 U5007 ( .B(\m5.addrM64 [61]), .A(n3432), .Z(n2306) );
  CANR1X1 U5008 ( .A(n3434), .B(\m0.addrM64 [61]), .C(n2306), .Z(n2307) );
  CND3X2 U5009 ( .A(n2309), .B(n2308), .C(n2307), .Z(n4151) );
  CAN2X1 U5010 ( .A(\s14.addr[18] ), .B(n4151), .Z(\s14.addr [61]) );
  CIVX2 U5011 ( .A(n2312), .Z(n2317) );
  CNR2X2 U5012 ( .A(n2314), .B(n2313), .Z(n2316) );
  CANR1X4 U5013 ( .A(n2317), .B(n2316), .C(n2315), .Z(n2318) );
  CIVX8 U5014 ( .A(n2318), .Z(n3417) );
  CIVX16 U5015 ( .A(n3417), .Z(\s11.en ) );
  CND2X1 U5016 ( .A(n3434), .B(\m0.addrM64 [29]), .Z(n2320) );
  CND2XL U5017 ( .A(n3436), .B(\m2.addrM64 [29]), .Z(n2319) );
  CND2X1 U5018 ( .A(n2320), .B(n2319), .Z(n2322) );
  CNR2X1 U5019 ( .A(n2322), .B(n2321), .Z(n2326) );
  CNR2IX1 U5020 ( .B(\m4.addrM64 [29]), .A(n3439), .Z(n2323) );
  CANR1X1 U5021 ( .A(n3431), .B(\m1.addrM64 [29]), .C(n2323), .Z(n2325) );
  CND2X1 U5022 ( .A(n3361), .B(\m3.addrM64 [29]), .Z(n2324) );
  CND3X2 U5023 ( .A(n2326), .B(n2325), .C(n2324), .Z(n4134) );
  CAN2XL U5024 ( .A(\s11.addr[17] ), .B(n4134), .Z(\s11.addr [29]) );
  CAN2XL U5025 ( .A(\s11.addr[17] ), .B(n4335), .Z(\s11.addr [8]) );
  CNR2IX1 U5026 ( .B(\m4.DoutM [23]), .A(n3439), .Z(n2327) );
  CNR2X1 U5027 ( .A(n2328), .B(n2327), .Z(n2333) );
  CANR2X1 U5028 ( .A(n3420), .B(\m3.DoutM [23]), .C(\m6.DoutM [23]), .D(n3435), 
        .Z(n2332) );
  CND2X1 U5029 ( .A(n3434), .B(\m0.DoutM [23]), .Z(n2330) );
  CNR2IX1 U5030 ( .B(\m5.DoutM [23]), .A(n3432), .Z(n2329) );
  CNR2IX1 U5031 ( .B(n2330), .A(n2329), .Z(n2331) );
  CND3X2 U5032 ( .A(n2333), .B(n2332), .C(n2331), .Z(n3483) );
  CAN2XL U5033 ( .A(\s11.addr[17] ), .B(n3483), .Z(\s11.SbusIn [23]) );
  CND2X1 U5034 ( .A(n3431), .B(\m1.DoutM [4]), .Z(n2335) );
  CND2XL U5035 ( .A(n3436), .B(\m2.DoutM [4]), .Z(n2334) );
  CND2X1 U5036 ( .A(n2335), .B(n2334), .Z(n2337) );
  CNR2IX1 U5037 ( .B(\m4.DoutM [4]), .A(n3439), .Z(n2336) );
  CNR2X1 U5038 ( .A(n2337), .B(n2336), .Z(n2341) );
  CANR2X1 U5039 ( .A(n3420), .B(\m3.DoutM [4]), .C(\m6.DoutM [4]), .D(n3435), 
        .Z(n2340) );
  CNR2IX1 U5040 ( .B(\m5.DoutM [4]), .A(n3432), .Z(n2338) );
  CANR1X1 U5041 ( .A(n3434), .B(\m0.DoutM [4]), .C(n2338), .Z(n2339) );
  CND3X2 U5042 ( .A(n2341), .B(n2340), .C(n2339), .Z(n4243) );
  CAN2X1 U5043 ( .A(\s7.en ), .B(n4243), .Z(\s7.SbusIn [4]) );
  CAN2X1 U5044 ( .A(\s7.en ), .B(n4180), .Z(\s7.SbusIn [18]) );
  CNIVX1 U5045 ( .A(n2342), .Z(n3289) );
  CND2X1 U5046 ( .A(n3289), .B(\m3.DoutM [19]), .Z(n2345) );
  CND2X1 U5047 ( .A(n3434), .B(\m0.DoutM [19]), .Z(n2344) );
  CND2X1 U5048 ( .A(n3431), .B(\m1.DoutM [19]), .Z(n2343) );
  CAN3X2 U5049 ( .A(n2345), .B(n2344), .C(n2343), .Z(n2353) );
  CIVX2 U5050 ( .A(\m5.DoutM [19]), .Z(n2347) );
  CND2X1 U5051 ( .A(n3435), .B(\m6.DoutM [19]), .Z(n2346) );
  CIVX2 U5052 ( .A(\m4.DoutM [19]), .Z(n2349) );
  CND2X1 U5053 ( .A(n3436), .B(\m2.DoutM [19]), .Z(n2348) );
  CNR2X1 U5054 ( .A(n2351), .B(n2350), .Z(n2352) );
  CND2X2 U5055 ( .A(n2353), .B(n2352), .Z(n4152) );
  CAN2X1 U5056 ( .A(\s7.addr[16] ), .B(n4152), .Z(\s7.SbusIn [19]) );
  CIVX8 U5057 ( .A(n3451), .Z(n4336) );
  CAN2X1 U5058 ( .A(n4336), .B(n3484), .Z(\s7.addr [11]) );
  CND2X1 U5059 ( .A(n3434), .B(\m0.DoutM [33]), .Z(n2355) );
  CND2XL U5060 ( .A(n3436), .B(\m2.DoutM [33]), .Z(n2354) );
  CND2X1 U5061 ( .A(n2355), .B(n2354), .Z(n2357) );
  CNR2X1 U5062 ( .A(n2357), .B(n2356), .Z(n2361) );
  CNR2IX1 U5063 ( .B(\m4.DoutM [33]), .A(n3439), .Z(n2358) );
  CANR1X1 U5064 ( .A(n3431), .B(\m1.DoutM [33]), .C(n2358), .Z(n2360) );
  CND2X1 U5065 ( .A(n3420), .B(\m3.DoutM [33]), .Z(n2359) );
  CND3X2 U5066 ( .A(n2361), .B(n2360), .C(n2359), .Z(n4156) );
  CAN2X1 U5067 ( .A(\s7.en ), .B(n4156), .Z(\s7.SbusIn [33]) );
  CND2X1 U5068 ( .A(n3289), .B(\m3.DoutM [25]), .Z(n2364) );
  CND2XL U5069 ( .A(n3434), .B(\m0.DoutM [25]), .Z(n2363) );
  CND2X1 U5070 ( .A(n3431), .B(\m1.DoutM [25]), .Z(n2362) );
  CAN3X2 U5071 ( .A(n2364), .B(n2363), .C(n2362), .Z(n2372) );
  CIVX2 U5072 ( .A(\m5.DoutM [25]), .Z(n2366) );
  CND2X1 U5073 ( .A(n3435), .B(\m6.DoutM [25]), .Z(n2365) );
  CIVX2 U5074 ( .A(\m4.DoutM [25]), .Z(n2368) );
  CND2X1 U5075 ( .A(n3436), .B(\m2.DoutM [25]), .Z(n2367) );
  CNR2X1 U5076 ( .A(n2370), .B(n2369), .Z(n2371) );
  CND2X2 U5077 ( .A(n2372), .B(n2371), .Z(n4141) );
  CAN2X1 U5078 ( .A(\s7.en ), .B(n4141), .Z(\s7.SbusIn [25]) );
  CNR2IX1 U5079 ( .B(\m5.DoutM [35]), .A(n3432), .Z(n2373) );
  CANR1X1 U5080 ( .A(n3431), .B(\m1.DoutM [35]), .C(n2373), .Z(n2378) );
  CNR2IX1 U5081 ( .B(\m4.DoutM [35]), .A(n3439), .Z(n2374) );
  CIVX2 U5082 ( .A(n2374), .Z(n2377) );
  CANR2X1 U5083 ( .A(n3435), .B(\m6.DoutM [35]), .C(\m3.DoutM [35]), .D(n3289), 
        .Z(n2376) );
  CANR2X1 U5084 ( .A(n3434), .B(\m0.DoutM [35]), .C(n3436), .D(\m2.DoutM [35]), 
        .Z(n2375) );
  CND4X4 U5085 ( .A(n2378), .B(n2377), .C(n2376), .D(n2375), .Z(n4237) );
  CAN2X1 U5086 ( .A(\s7.addr[16] ), .B(n4237), .Z(\s7.SbusIn [35]) );
  CAN2X1 U5087 ( .A(n4336), .B(n4121), .Z(\s7.SbusIn [48]) );
  CND2X1 U5088 ( .A(n3431), .B(\m1.DoutM [39]), .Z(n2380) );
  CND2XL U5089 ( .A(n3436), .B(\m2.DoutM [39]), .Z(n2379) );
  CND2X1 U5090 ( .A(n2380), .B(n2379), .Z(n2382) );
  CNR2IX1 U5091 ( .B(\m4.DoutM [39]), .A(n3439), .Z(n2381) );
  CNR2X1 U5092 ( .A(n2382), .B(n2381), .Z(n2386) );
  CANR2X1 U5093 ( .A(n1842), .B(\m3.DoutM [39]), .C(\m6.DoutM [39]), .D(n3435), 
        .Z(n2385) );
  CNR2IX1 U5094 ( .B(\m5.DoutM [39]), .A(n3432), .Z(n2383) );
  CANR1X1 U5095 ( .A(n3434), .B(\m0.DoutM [39]), .C(n2383), .Z(n2384) );
  CND3X2 U5096 ( .A(n2386), .B(n2385), .C(n2384), .Z(n4135) );
  CAN2X1 U5097 ( .A(\s7.en ), .B(n4135), .Z(\s7.SbusIn [39]) );
  CND2X1 U5098 ( .A(n3434), .B(\m0.DoutM [30]), .Z(n2388) );
  CND2X1 U5099 ( .A(n3436), .B(\m2.DoutM [30]), .Z(n2387) );
  CND2X1 U5100 ( .A(n2388), .B(n2387), .Z(n2392) );
  CIVX2 U5101 ( .A(\m5.DoutM [30]), .Z(n2390) );
  CND2X1 U5102 ( .A(n3435), .B(\m6.DoutM [30]), .Z(n2389) );
  CNR2X1 U5103 ( .A(n2392), .B(n2391), .Z(n2396) );
  CANR2X1 U5104 ( .A(n3431), .B(\m1.DoutM [30]), .C(\m3.DoutM [30]), .D(n3137), 
        .Z(n2395) );
  CNR2IX1 U5105 ( .B(\m4.DoutM [30]), .A(n3439), .Z(n2393) );
  CIVX2 U5106 ( .A(n2393), .Z(n2394) );
  CAN2X1 U5107 ( .A(\s7.addr[19] ), .B(n4145), .Z(\s7.SbusIn [30]) );
  CANR2X1 U5108 ( .A(n3431), .B(\m1.DoutM [20]), .C(\m3.DoutM [20]), .D(n3137), 
        .Z(n2404) );
  CNR2IX1 U5109 ( .B(\m5.DoutM [20]), .A(n3432), .Z(n2397) );
  CANR1X1 U5110 ( .A(n3434), .B(\m0.DoutM [20]), .C(n2397), .Z(n2403) );
  CND2XL U5111 ( .A(n3435), .B(\m6.DoutM [20]), .Z(n2399) );
  CND2X1 U5112 ( .A(n3436), .B(\m2.DoutM [20]), .Z(n2398) );
  CND2X1 U5113 ( .A(n2399), .B(n2398), .Z(n2401) );
  CNR2IX1 U5114 ( .B(\m4.DoutM [20]), .A(n3439), .Z(n2400) );
  CNR2X2 U5115 ( .A(n2401), .B(n2400), .Z(n2402) );
  CND3X2 U5116 ( .A(n2404), .B(n2403), .C(n2402), .Z(n4150) );
  CAN2X1 U5117 ( .A(\s7.addr[16] ), .B(n4150), .Z(\s7.SbusIn [20]) );
  CND2XL U5118 ( .A(n3431), .B(\m1.DoutM [13]), .Z(n2406) );
  CND2XL U5119 ( .A(n3436), .B(\m2.DoutM [13]), .Z(n2405) );
  CND2X1 U5120 ( .A(n2406), .B(n2405), .Z(n2408) );
  CNR2IX1 U5121 ( .B(\m4.DoutM [13]), .A(n3439), .Z(n2407) );
  CNR2X1 U5122 ( .A(n2408), .B(n2407), .Z(n2412) );
  CANR2X1 U5123 ( .A(n3299), .B(\m3.DoutM [13]), .C(\m6.DoutM [13]), .D(n3435), 
        .Z(n2411) );
  CNR2IX1 U5124 ( .B(\m5.DoutM [13]), .A(n3432), .Z(n2409) );
  CANR1X1 U5125 ( .A(n3434), .B(\m0.DoutM [13]), .C(n2409), .Z(n2410) );
  CND3X2 U5126 ( .A(n2412), .B(n2411), .C(n2410), .Z(n4123) );
  CAN2X1 U5127 ( .A(n4336), .B(n4123), .Z(\s7.SbusIn [13]) );
  CNR2IX1 U5128 ( .B(\m4.DoutM [46]), .A(n3439), .Z(n2413) );
  CNR2X1 U5129 ( .A(n2414), .B(n2413), .Z(n2418) );
  CANR2X1 U5130 ( .A(n3435), .B(\m6.DoutM [46]), .C(\m3.DoutM [46]), .D(n3361), 
        .Z(n2417) );
  CNR2IX1 U5131 ( .B(\m5.DoutM [46]), .A(n3432), .Z(n2415) );
  CND3X2 U5132 ( .A(n2418), .B(n2417), .C(n2416), .Z(n3472) );
  CAN2X1 U5133 ( .A(\s7.addr[19] ), .B(n3472), .Z(\s7.SbusIn [46]) );
  CND2X1 U5134 ( .A(n3431), .B(\m1.DoutM [53]), .Z(n2420) );
  CND2XL U5135 ( .A(n3436), .B(\m2.DoutM [53]), .Z(n2419) );
  CND2X1 U5136 ( .A(n2420), .B(n2419), .Z(n2422) );
  CNR2IX1 U5137 ( .B(\m4.DoutM [53]), .A(n3439), .Z(n2421) );
  CNR2X1 U5138 ( .A(n2422), .B(n2421), .Z(n2426) );
  CANR2X1 U5139 ( .A(n3361), .B(\m3.DoutM [53]), .C(\m6.DoutM [53]), .D(n3435), 
        .Z(n2425) );
  CNR2IX1 U5140 ( .B(\m5.DoutM [53]), .A(n3432), .Z(n2423) );
  CND3X2 U5141 ( .A(n2426), .B(n2425), .C(n2424), .Z(n4170) );
  CAN2X1 U5142 ( .A(\s7.en ), .B(n4170), .Z(\s7.SbusIn [53]) );
  CAN2X1 U5143 ( .A(\s7.addr[16] ), .B(n4335), .Z(\s7.addr [8]) );
  CANR2X1 U5144 ( .A(n3431), .B(\m1.DoutM [1]), .C(\m3.DoutM [1]), .D(n3420), 
        .Z(n2434) );
  CNR2IX1 U5145 ( .B(\m5.DoutM [1]), .A(n3432), .Z(n2427) );
  CANR1X1 U5146 ( .A(n3434), .B(\m0.DoutM [1]), .C(n2427), .Z(n2433) );
  CND2X1 U5147 ( .A(n3435), .B(\m6.DoutM [1]), .Z(n2429) );
  CND2X1 U5148 ( .A(n3436), .B(\m2.DoutM [1]), .Z(n2428) );
  CND2X1 U5149 ( .A(n2429), .B(n2428), .Z(n2431) );
  CNR2IX1 U5150 ( .B(\m4.DoutM [1]), .A(n3439), .Z(n2430) );
  CNR2X1 U5151 ( .A(n2431), .B(n2430), .Z(n2432) );
  CND3X2 U5152 ( .A(n2434), .B(n2433), .C(n2432), .Z(n4190) );
  CAN2X1 U5153 ( .A(\s7.addr[19] ), .B(n4190), .Z(\s7.SbusIn [1]) );
  CIVX20 U5154 ( .A(n3415), .Z(\s8.addr[17] ) );
  CNR2IX1 U5155 ( .B(\m5.DoutM [7]), .A(n3432), .Z(n2436) );
  CNR2IX1 U5156 ( .B(\m4.DoutM [7]), .A(n3439), .Z(n2437) );
  CIVX2 U5157 ( .A(n2437), .Z(n2441) );
  CANR2X1 U5158 ( .A(n3435), .B(\m6.DoutM [7]), .C(\m3.DoutM [7]), .D(n3371), 
        .Z(n2440) );
  CAN2X1 U5159 ( .A(n3436), .B(\m2.DoutM [7]), .Z(n2438) );
  CND4X2 U5160 ( .A(n2442), .B(n2441), .C(n2440), .D(n2439), .Z(n4154) );
  CAN2X1 U5161 ( .A(\s8.addr[17] ), .B(n4154), .Z(\s8.SbusIn [7]) );
  CNR2IX1 U5162 ( .B(\m4.DoutM [2]), .A(n3439), .Z(n2443) );
  CNR2X1 U5163 ( .A(n2444), .B(n2443), .Z(n2449) );
  CANR2X1 U5164 ( .A(n3430), .B(\m3.DoutM [2]), .C(\m6.DoutM [2]), .D(n3435), 
        .Z(n2448) );
  CND2X1 U5165 ( .A(n3434), .B(\m0.DoutM [2]), .Z(n2446) );
  CNR2IX1 U5166 ( .B(\m5.DoutM [2]), .A(n3432), .Z(n2445) );
  CNR2IX1 U5167 ( .B(n2446), .A(n2445), .Z(n2447) );
  CND3X2 U5168 ( .A(n2449), .B(n2448), .C(n2447), .Z(n4192) );
  CAN2XL U5169 ( .A(\s6.en ), .B(n4192), .Z(\s6.SbusIn [2]) );
  CIVX2 U5170 ( .A(n2452), .Z(n2453) );
  CND2X4 U5171 ( .A(n2454), .B(n2453), .Z(n2455) );
  COND4CX1 U5172 ( .A(n3468), .B(n2754), .C(n2780), .D(n2789), .Z(n2457) );
  CAN2X1 U5173 ( .A(n3454), .B(n2459), .Z(n2460) );
  CAN2X2 U5174 ( .A(n2461), .B(n2460), .Z(n2468) );
  CNR2X2 U5175 ( .A(n2462), .B(n2731), .Z(n2463) );
  CND3X2 U5176 ( .A(n2465), .B(n2464), .C(n2463), .Z(n2466) );
  CIVX4 U5177 ( .A(n2466), .Z(n2760) );
  CND3X4 U5178 ( .A(n2468), .B(n2760), .C(n2467), .Z(n2469) );
  CIVX8 U5179 ( .A(n2469), .Z(n2511) );
  CND2X4 U5180 ( .A(n2512), .B(n2511), .Z(n2812) );
  CIVDX2 U5181 ( .A(n2470), .Z0(n2139), .Z1(n3485) );
  CAN2X1 U5182 ( .A(n4405), .B(n3485), .Z(\s5.addr [6]) );
  CAN2X1 U5183 ( .A(n1844), .B(n4156), .Z(\s5.SbusIn [33]) );
  CND2X1 U5184 ( .A(n3434), .B(\m0.DoutM [51]), .Z(n2472) );
  CND2X1 U5185 ( .A(n3436), .B(\m2.DoutM [51]), .Z(n2471) );
  CND2X1 U5186 ( .A(n2472), .B(n2471), .Z(n2474) );
  CNR2X1 U5187 ( .A(n2474), .B(n2473), .Z(n2478) );
  CNR2IX1 U5188 ( .B(\m4.DoutM [51]), .A(n3439), .Z(n2475) );
  CANR1X1 U5189 ( .A(n3431), .B(\m1.DoutM [51]), .C(n2475), .Z(n2477) );
  CND2X1 U5190 ( .A(n3137), .B(\m3.DoutM [51]), .Z(n2476) );
  CND3X2 U5191 ( .A(n2478), .B(n2477), .C(n2476), .Z(n4163) );
  CAN2X1 U5192 ( .A(n5445), .B(n4163), .Z(\s5.SbusIn [51]) );
  CANR2X1 U5193 ( .A(n3431), .B(\m1.addrM64 [48]), .C(\m3.addrM64 [48]), .D(
        n3420), .Z(n2486) );
  CNR2IX1 U5194 ( .B(\m5.addrM64 [48]), .A(n3432), .Z(n2479) );
  CANR1X1 U5195 ( .A(n3434), .B(\m0.addrM64 [48]), .C(n2479), .Z(n2485) );
  CND2XL U5196 ( .A(n3435), .B(\m6.addrM64 [48]), .Z(n2481) );
  CND2X1 U5197 ( .A(n3436), .B(\m2.addrM64 [48]), .Z(n2480) );
  CND2X1 U5198 ( .A(n2481), .B(n2480), .Z(n2483) );
  CNR2IX1 U5199 ( .B(\m4.addrM64 [48]), .A(n3439), .Z(n2482) );
  CNR2X2 U5200 ( .A(n2483), .B(n2482), .Z(n2484) );
  CND3X2 U5201 ( .A(n2486), .B(n2485), .C(n2484), .Z(n4137) );
  CAN2X1 U5202 ( .A(n4405), .B(n4137), .Z(\s5.addr [48]) );
  CAN2X1 U5203 ( .A(n4405), .B(n4170), .Z(\s5.SbusIn [53]) );
  CND2X1 U5204 ( .A(n3434), .B(\m0.addrM64 [20]), .Z(n2488) );
  CND2XL U5205 ( .A(n3436), .B(\m2.addrM64 [20]), .Z(n2487) );
  CND2X1 U5206 ( .A(n2488), .B(n2487), .Z(n2490) );
  CNR2X1 U5207 ( .A(n2490), .B(n2489), .Z(n2494) );
  CNR2IX1 U5208 ( .B(\m4.addrM64 [20]), .A(n3439), .Z(n2491) );
  CANR1X1 U5209 ( .A(n3431), .B(\m1.addrM64 [20]), .C(n2491), .Z(n2493) );
  CND2X1 U5210 ( .A(n3420), .B(\m3.addrM64 [20]), .Z(n2492) );
  CND3X2 U5211 ( .A(n2494), .B(n2493), .C(n2492), .Z(n4331) );
  CAN2X1 U5212 ( .A(n4405), .B(n4331), .Z(\s5.addr [20]) );
  CND2XL U5213 ( .A(n3431), .B(\m1.DoutM [59]), .Z(n2496) );
  CND2XL U5214 ( .A(n3436), .B(\m2.DoutM [59]), .Z(n2495) );
  CND2X1 U5215 ( .A(n2496), .B(n2495), .Z(n2498) );
  CNR2IX1 U5216 ( .B(\m4.DoutM [59]), .A(n3439), .Z(n2497) );
  CNR2X1 U5217 ( .A(n2498), .B(n2497), .Z(n2502) );
  CANR2X1 U5218 ( .A(n3289), .B(\m3.DoutM [59]), .C(\m6.DoutM [59]), .D(n3435), 
        .Z(n2501) );
  CNR2IX1 U5219 ( .B(\m5.DoutM [59]), .A(n3432), .Z(n2499) );
  CND3X2 U5220 ( .A(n2502), .B(n2501), .C(n2500), .Z(n4130) );
  CAN2X1 U5221 ( .A(n4405), .B(n4130), .Z(\s5.SbusIn [59]) );
  CANR2X1 U5222 ( .A(n3431), .B(\m1.DoutM [62]), .C(\m3.DoutM [62]), .D(n3289), 
        .Z(n2510) );
  CNR2IX1 U5223 ( .B(\m5.DoutM [62]), .A(n3432), .Z(n2503) );
  CANR1X1 U5224 ( .A(n3434), .B(\m0.DoutM [62]), .C(n2503), .Z(n2509) );
  CND2XL U5225 ( .A(n3435), .B(\m6.DoutM [62]), .Z(n2505) );
  CND2X1 U5226 ( .A(n3436), .B(\m2.DoutM [62]), .Z(n2504) );
  CND2X1 U5227 ( .A(n2505), .B(n2504), .Z(n2507) );
  CNR2IX1 U5228 ( .B(\m4.DoutM [62]), .A(n3439), .Z(n2506) );
  CNR2X2 U5229 ( .A(n2507), .B(n2506), .Z(n2508) );
  CND3X2 U5230 ( .A(n2510), .B(n2509), .C(n2508), .Z(n4126) );
  CAN2X1 U5231 ( .A(n1844), .B(n4126), .Z(\s5.SbusIn [62]) );
  CND2X4 U5232 ( .A(n2512), .B(n2511), .Z(n2513) );
  CND2X1 U5233 ( .A(n3431), .B(\m1.DoutM [44]), .Z(n2515) );
  CND2XL U5234 ( .A(n3436), .B(\m2.DoutM [44]), .Z(n2514) );
  CND2X1 U5235 ( .A(n2515), .B(n2514), .Z(n2517) );
  CNR2IX1 U5236 ( .B(\m4.DoutM [44]), .A(n3439), .Z(n2516) );
  CNR2X1 U5237 ( .A(n2517), .B(n2516), .Z(n2521) );
  CANR2X1 U5238 ( .A(n3289), .B(\m3.DoutM [44]), .C(\m6.DoutM [44]), .D(n3435), 
        .Z(n2520) );
  CNR2IX1 U5239 ( .B(\m5.DoutM [44]), .A(n3432), .Z(n2518) );
  CND3X2 U5240 ( .A(n2521), .B(n2520), .C(n2519), .Z(n4138) );
  CAN2X1 U5241 ( .A(n4405), .B(n4138), .Z(\s5.SbusIn [44]) );
  COND1X2 U5242 ( .A(n2790), .B(n2522), .C(n4257), .Z(n2526) );
  CND2X2 U5243 ( .A(n2523), .B(n2774), .Z(n2524) );
  CND2X4 U5244 ( .A(n3459), .B(n2524), .Z(n2751) );
  CIVX2 U5245 ( .A(n2751), .Z(n2545) );
  CND2X2 U5246 ( .A(n2789), .B(n2623), .Z(n2630) );
  CND3X2 U5247 ( .A(n2526), .B(n2525), .C(n2630), .Z(n2534) );
  CND3X1 U5248 ( .A(n2527), .B(n2761), .C(n5518), .Z(n2530) );
  CNR3X2 U5249 ( .A(n2530), .B(n2529), .C(n2528), .Z(n2531) );
  CND2X2 U5250 ( .A(n2760), .B(n2531), .Z(n2532) );
  CIVX2 U5251 ( .A(n2532), .Z(n2533) );
  CND2X4 U5252 ( .A(n2534), .B(n2533), .Z(n2535) );
  CIVX8 U5253 ( .A(n2535), .Z(n2536) );
  CIVX16 U5254 ( .A(n2536), .Z(n3445) );
  CIVX12 U5255 ( .A(n3445), .Z(\s4.addr[14] ) );
  CIVX16 U5256 ( .A(n3445), .Z(\s4.en ) );
  CAN2X2 U5257 ( .A(n2537), .B(n2548), .Z(n2540) );
  CNR2X2 U5258 ( .A(n2538), .B(n2645), .Z(n2539) );
  CNR2X4 U5259 ( .A(n2540), .B(n2539), .Z(n2808) );
  CND3X1 U5260 ( .A(n2543), .B(n2542), .C(n2541), .Z(n2544) );
  CNR2X2 U5261 ( .A(n2645), .B(n2544), .Z(n2546) );
  CND2X2 U5262 ( .A(n2546), .B(n2545), .Z(n2550) );
  CND3X2 U5263 ( .A(n2548), .B(n2547), .C(n2790), .Z(n2549) );
  CND2X2 U5264 ( .A(n2550), .B(n2549), .Z(n2551) );
  CIVX4 U5265 ( .A(n2551), .Z(n2809) );
  CNR2X2 U5266 ( .A(n2614), .B(\c1.Breset ), .Z(n2554) );
  CND2X2 U5267 ( .A(n2552), .B(n2729), .Z(n2612) );
  CNR2X4 U5268 ( .A(n2786), .B(n2612), .Z(n2553) );
  CND2X4 U5269 ( .A(n2554), .B(n2553), .Z(n2807) );
  CANR1X4 U5270 ( .A(n2808), .B(n2809), .C(n2807), .Z(n2555) );
  CIVX8 U5271 ( .A(n2555), .Z(n3416) );
  CIVX16 U5272 ( .A(n3416), .Z(\s10.addr[9] ) );
  CNR2IX1 U5273 ( .B(\m5.DoutM [26]), .A(n3432), .Z(n2556) );
  CNR2IX1 U5274 ( .B(\m4.DoutM [26]), .A(n3439), .Z(n2557) );
  CIVX2 U5275 ( .A(n2557), .Z(n2560) );
  CANR2X1 U5276 ( .A(n3361), .B(\m3.DoutM [26]), .C(\m6.DoutM [26]), .D(n3435), 
        .Z(n2559) );
  CANR2X1 U5277 ( .A(n3434), .B(\m0.DoutM [26]), .C(n3436), .D(\m2.DoutM [26]), 
        .Z(n2558) );
  CND4X2 U5278 ( .A(n2561), .B(n2560), .C(n2559), .D(n2558), .Z(n4147) );
  CAN2X1 U5279 ( .A(\s10.addr[9] ), .B(n4147), .Z(\s10.SbusIn [26]) );
  CND2X1 U5280 ( .A(n3431), .B(\m1.addrM64 [21]), .Z(n2563) );
  CND2XL U5281 ( .A(n3436), .B(\m2.addrM64 [21]), .Z(n2562) );
  CND2X1 U5282 ( .A(n2563), .B(n2562), .Z(n2565) );
  CNR2IX1 U5283 ( .B(\m4.addrM64 [21]), .A(n3439), .Z(n2564) );
  CNR2X1 U5284 ( .A(n2565), .B(n2564), .Z(n2569) );
  CANR2X1 U5285 ( .A(n3435), .B(\m6.addrM64 [21]), .C(\m3.addrM64 [21]), .D(
        n3420), .Z(n2568) );
  CNR2IX1 U5286 ( .B(\m5.addrM64 [21]), .A(n3432), .Z(n2566) );
  CND3X2 U5287 ( .A(n2569), .B(n2568), .C(n2567), .Z(n4128) );
  CAN2X1 U5288 ( .A(\s10.addr[9] ), .B(n4128), .Z(\s10.addr [21]) );
  CANR1X4 U5289 ( .A(n2808), .B(n2809), .C(n2807), .Z(n2570) );
  CIVX8 U5290 ( .A(n2570), .Z(n2571) );
  CIVX16 U5291 ( .A(n2571), .Z(\s10.en ) );
  CANR2X1 U5292 ( .A(n3431), .B(\m1.DoutM [12]), .C(\m3.DoutM [12]), .D(n3420), 
        .Z(n2579) );
  CNR2IX1 U5293 ( .B(\m5.DoutM [12]), .A(n3432), .Z(n2572) );
  CANR1X1 U5294 ( .A(n3434), .B(\m0.DoutM [12]), .C(n2572), .Z(n2578) );
  CND2X1 U5295 ( .A(n3435), .B(\m6.DoutM [12]), .Z(n2574) );
  CND2X1 U5296 ( .A(n3436), .B(\m2.DoutM [12]), .Z(n2573) );
  CND2X1 U5297 ( .A(n2574), .B(n2573), .Z(n2576) );
  CNR2IX1 U5298 ( .B(\m4.DoutM [12]), .A(n3439), .Z(n2575) );
  CNR2X1 U5299 ( .A(n2576), .B(n2575), .Z(n2577) );
  CND3X2 U5300 ( .A(n2579), .B(n2578), .C(n2577), .Z(n3481) );
  CAN2X1 U5301 ( .A(\s10.en ), .B(n3481), .Z(\s10.SbusIn [12]) );
  CND2X1 U5302 ( .A(n3434), .B(\m0.DoutM [0]), .Z(n2581) );
  CND2XL U5303 ( .A(n3436), .B(\m2.DoutM [0]), .Z(n2580) );
  CIVX2 U5304 ( .A(\m5.DoutM [0]), .Z(n2583) );
  CND2X1 U5305 ( .A(n3435), .B(\m6.DoutM [0]), .Z(n2582) );
  CAN2XL U5306 ( .A(\s10.en ), .B(n4185), .Z(\s10.SbusIn [0]) );
  CAN2XL U5307 ( .A(\s10.en ), .B(n4200), .Z(\s10.SbusIn [3]) );
  CAN2XL U5308 ( .A(\s10.en ), .B(n4135), .Z(\s10.SbusIn [39]) );
  CND2X1 U5309 ( .A(n3431), .B(\m1.DoutM [28]), .Z(n2585) );
  CND2XL U5310 ( .A(n3436), .B(\m2.DoutM [28]), .Z(n2584) );
  CND2X1 U5311 ( .A(n2585), .B(n2584), .Z(n2587) );
  CNR2IX1 U5312 ( .B(\m4.DoutM [28]), .A(n3439), .Z(n2586) );
  CNR2X1 U5313 ( .A(n2587), .B(n2586), .Z(n2591) );
  CANR2X1 U5314 ( .A(n3371), .B(\m3.DoutM [28]), .C(\m6.DoutM [28]), .D(n3435), 
        .Z(n2590) );
  CNR2IX1 U5315 ( .B(\m5.DoutM [28]), .A(n3432), .Z(n2588) );
  CANR1X1 U5316 ( .A(n3434), .B(\m0.DoutM [28]), .C(n2588), .Z(n2589) );
  CND3X2 U5317 ( .A(n2591), .B(n2590), .C(n2589), .Z(n4117) );
  CAN2XL U5318 ( .A(\s10.en ), .B(n4117), .Z(\s10.SbusIn [28]) );
  CND2X1 U5319 ( .A(n3434), .B(\m0.DoutM [32]), .Z(n2593) );
  CND2XL U5320 ( .A(n3436), .B(\m2.DoutM [32]), .Z(n2592) );
  CND2X1 U5321 ( .A(n2593), .B(n2592), .Z(n2597) );
  CIVX2 U5322 ( .A(\m5.DoutM [32]), .Z(n2595) );
  CND2X1 U5323 ( .A(n3435), .B(\m6.DoutM [32]), .Z(n2594) );
  CNR2X1 U5324 ( .A(n2597), .B(n2596), .Z(n2601) );
  CANR2X1 U5325 ( .A(n3431), .B(\m1.DoutM [32]), .C(\m3.DoutM [32]), .D(n3420), 
        .Z(n2600) );
  CNR2IX1 U5326 ( .B(\m4.DoutM [32]), .A(n3439), .Z(n2598) );
  CIVX2 U5327 ( .A(n2598), .Z(n2599) );
  CAN2XL U5328 ( .A(\s10.en ), .B(n4171), .Z(\s10.SbusIn [32]) );
  CND2X1 U5329 ( .A(n3434), .B(\m0.DoutM [34]), .Z(n2603) );
  CND2XL U5330 ( .A(n3436), .B(\m2.DoutM [34]), .Z(n2602) );
  CND2X1 U5331 ( .A(n2603), .B(n2602), .Z(n2607) );
  CIVX2 U5332 ( .A(\m5.DoutM [34]), .Z(n2605) );
  CND2X1 U5333 ( .A(n3435), .B(\m6.DoutM [34]), .Z(n2604) );
  CNR2X1 U5334 ( .A(n2607), .B(n2606), .Z(n2611) );
  CANR2X1 U5335 ( .A(n3431), .B(\m1.DoutM [34]), .C(\m3.DoutM [34]), .D(n3289), 
        .Z(n2610) );
  CNR2IX1 U5336 ( .B(\m4.DoutM [34]), .A(n3439), .Z(n2608) );
  CIVX2 U5337 ( .A(n2608), .Z(n2609) );
  CAN2XL U5338 ( .A(\s10.en ), .B(n4178), .Z(\s10.SbusIn [34]) );
  CNR2X2 U5339 ( .A(n2786), .B(n2612), .Z(n2617) );
  CNR2IX2 U5340 ( .B(n2615), .A(n2614), .Z(n2616) );
  CND3X2 U5341 ( .A(n2618), .B(n2617), .C(n2616), .Z(n2619) );
  CIVX2 U5342 ( .A(n2619), .Z(n2627) );
  COND1X1 U5343 ( .A(n2751), .B(n2620), .C(n2789), .Z(n2625) );
  CND4X1 U5344 ( .A(n2793), .B(n2623), .C(n2622), .D(n2621), .Z(n2624) );
  CND2X2 U5345 ( .A(n2625), .B(n2624), .Z(n2626) );
  CND2X4 U5346 ( .A(n2627), .B(n2626), .Z(n2628) );
  CIVX12 U5347 ( .A(n2628), .Z(n3463) );
  CIVX20 U5348 ( .A(n3463), .Z(n3298) );
  CIVX20 U5349 ( .A(n3298), .Z(\s9.addr[8] ) );
  CNR2X2 U5350 ( .A(n2630), .B(n2629), .Z(n2644) );
  CIVDX2 U5351 ( .A(n2631), .Z0(n4326), .Z1(n3478) );
  CND3X4 U5352 ( .A(n2638), .B(n2637), .C(n2636), .Z(n4330) );
  CIVX8 U5353 ( .A(n4330), .Z(n4318) );
  CND2X4 U5354 ( .A(n4318), .B(n3459), .Z(n2640) );
  CND3X4 U5355 ( .A(n2640), .B(n3476), .C(n2639), .Z(n2641) );
  CANR1X4 U5356 ( .A(n2642), .B(n2641), .C(n3456), .Z(n2643) );
  CNR2X4 U5357 ( .A(n2644), .B(n2643), .Z(n2721) );
  CIVX2 U5358 ( .A(n2721), .Z(n2649) );
  CNR2IX1 U5359 ( .B(n5518), .A(n2645), .Z(n2646) );
  CND2X2 U5360 ( .A(n2647), .B(n2646), .Z(n2720) );
  CIVX2 U5361 ( .A(n2720), .Z(n2648) );
  CND2X4 U5362 ( .A(n2649), .B(n2648), .Z(n3446) );
  CIVX16 U5363 ( .A(n3446), .Z(\s1.addr[17] ) );
  CND2X1 U5364 ( .A(n3434), .B(\m0.DoutM [11]), .Z(n2651) );
  CND2XL U5365 ( .A(n3436), .B(\m2.DoutM [11]), .Z(n2650) );
  CND2X1 U5366 ( .A(n2651), .B(n2650), .Z(n2653) );
  CNR2X1 U5367 ( .A(n2653), .B(n2652), .Z(n2657) );
  CNR2IX1 U5368 ( .B(\m4.DoutM [11]), .A(n3439), .Z(n2654) );
  CANR1X1 U5369 ( .A(n3431), .B(\m1.DoutM [11]), .C(n2654), .Z(n2656) );
  CND2X1 U5370 ( .A(n3371), .B(\m3.DoutM [11]), .Z(n2655) );
  CND3X2 U5371 ( .A(n2657), .B(n2656), .C(n2655), .Z(n3465) );
  CAN2XL U5372 ( .A(\s6.addr [17]), .B(n3465), .Z(\s6.SbusIn [11]) );
  CAN2XL U5373 ( .A(\s6.addr [17]), .B(n4243), .Z(\s6.SbusIn [4]) );
  CNR2IX1 U5374 ( .B(\m5.addrM64 [56]), .A(n3432), .Z(n2658) );
  CND2XL U5375 ( .A(n3424), .B(\m4.addrM64 [56]), .Z(n2661) );
  CANR2X1 U5376 ( .A(n3371), .B(\m3.addrM64 [56]), .C(\m6.addrM64 [56]), .D(
        n3435), .Z(n2660) );
  CANR2X1 U5377 ( .A(n3434), .B(\m0.addrM64 [56]), .C(n3436), .D(
        \m2.addrM64 [56]), .Z(n2659) );
  CND4X2 U5378 ( .A(n2662), .B(n2661), .C(n2660), .D(n2659), .Z(n4242) );
  CAN2XL U5379 ( .A(\s6.addr [17]), .B(n4242), .Z(\s6.addr [56]) );
  CND2XL U5380 ( .A(n3361), .B(\m3.addrM64 [55]), .Z(n2665) );
  CND2X1 U5381 ( .A(n3434), .B(\m0.addrM64 [55]), .Z(n2664) );
  CND2X1 U5382 ( .A(n3431), .B(\m1.addrM64 [55]), .Z(n2663) );
  CAN3X2 U5383 ( .A(n2665), .B(n2664), .C(n2663), .Z(n2673) );
  CIVX2 U5384 ( .A(\m5.addrM64 [55]), .Z(n2667) );
  CND2X1 U5385 ( .A(n3435), .B(\m6.addrM64 [55]), .Z(n2666) );
  CIVX2 U5386 ( .A(\m4.addrM64 [55]), .Z(n2669) );
  CND2X1 U5387 ( .A(n3436), .B(\m2.addrM64 [55]), .Z(n2668) );
  CNR2X1 U5388 ( .A(n2671), .B(n2670), .Z(n2672) );
  CND2X2 U5389 ( .A(n2673), .B(n2672), .Z(n4201) );
  CAN2XL U5390 ( .A(\s6.addr [17]), .B(n4201), .Z(\s6.addr [55]) );
  CND2XL U5391 ( .A(n2855), .B(\m3.DoutM [61]), .Z(n2676) );
  CND2X1 U5392 ( .A(n3434), .B(\m0.DoutM [61]), .Z(n2675) );
  CND2X1 U5393 ( .A(n3431), .B(\m1.DoutM [61]), .Z(n2674) );
  CAN3X2 U5394 ( .A(n2676), .B(n2675), .C(n2674), .Z(n2682) );
  CIVX2 U5395 ( .A(\m5.DoutM [61]), .Z(n2678) );
  CND2X1 U5396 ( .A(n3435), .B(\m6.DoutM [61]), .Z(n2677) );
  CNR2X1 U5397 ( .A(n2680), .B(n2679), .Z(n2681) );
  CND2X2 U5398 ( .A(n2682), .B(n2681), .Z(n4125) );
  CAN2XL U5399 ( .A(\s6.addr [17]), .B(n4125), .Z(\s6.SbusIn [61]) );
  CIVX2 U5400 ( .A(\m5.DoutM [60]), .Z(n2684) );
  CND2X1 U5401 ( .A(n3435), .B(\m6.DoutM [60]), .Z(n2683) );
  COND1X1 U5402 ( .A(n3432), .B(n2684), .C(n2683), .Z(n2685) );
  CNR2X1 U5403 ( .A(n2686), .B(n2685), .Z(n2690) );
  CNR2IX1 U5404 ( .B(\m4.DoutM [60]), .A(n3439), .Z(n2687) );
  CANR1X1 U5405 ( .A(n3431), .B(\m1.DoutM [60]), .C(n2687), .Z(n2689) );
  CND2X1 U5406 ( .A(n3420), .B(\m3.DoutM [60]), .Z(n2688) );
  CND3X2 U5407 ( .A(n2690), .B(n2689), .C(n2688), .Z(n4167) );
  CAN2XL U5408 ( .A(\s6.addr [17]), .B(n4167), .Z(\s6.SbusIn [60]) );
  CAN2XL U5409 ( .A(\s6.addr [17]), .B(n4163), .Z(\s6.SbusIn [51]) );
  CANR2X1 U5410 ( .A(n3431), .B(\m1.DoutM [50]), .C(\m3.DoutM [50]), .D(n3371), 
        .Z(n2698) );
  CNR2IX1 U5411 ( .B(\m5.DoutM [50]), .A(n3432), .Z(n2691) );
  CANR1X1 U5412 ( .A(n3434), .B(\m0.DoutM [50]), .C(n2691), .Z(n2697) );
  CND2XL U5413 ( .A(n3435), .B(\m6.DoutM [50]), .Z(n2693) );
  CND2X1 U5414 ( .A(n3436), .B(\m2.DoutM [50]), .Z(n2692) );
  CND2X1 U5415 ( .A(n2693), .B(n2692), .Z(n2695) );
  CNR2IX1 U5416 ( .B(\m4.DoutM [50]), .A(n3439), .Z(n2694) );
  CNR2X1 U5417 ( .A(n2695), .B(n2694), .Z(n2696) );
  CND3X2 U5418 ( .A(n2698), .B(n2697), .C(n2696), .Z(n4127) );
  CAN2XL U5419 ( .A(\s6.addr [17]), .B(n4127), .Z(\s6.SbusIn [50]) );
  CANR2X1 U5420 ( .A(n3431), .B(\m1.DoutM [22]), .C(\m3.DoutM [22]), .D(n3299), 
        .Z(n2705) );
  CND2X1 U5421 ( .A(n3434), .B(\m0.DoutM [22]), .Z(n2700) );
  CNR2IX1 U5422 ( .B(\m5.DoutM [22]), .A(n3432), .Z(n2699) );
  CNR2IX1 U5423 ( .B(n2700), .A(n2699), .Z(n2704) );
  CNR2IX1 U5424 ( .B(\m4.DoutM [22]), .A(n3439), .Z(n2701) );
  CNR2X1 U5425 ( .A(n2702), .B(n2701), .Z(n2703) );
  CND3X2 U5426 ( .A(n2705), .B(n2704), .C(n2703), .Z(n3473) );
  CAN2XL U5427 ( .A(\s6.addr [17]), .B(n3473), .Z(\s6.SbusIn [22]) );
  CAN2XL U5428 ( .A(\s6.addr [17]), .B(n4150), .Z(\s6.SbusIn [20]) );
  CNR2IX1 U5429 ( .B(\m5.addrM64 [36]), .A(n3432), .Z(n2706) );
  CNR2IX1 U5430 ( .B(\m4.addrM64 [36]), .A(n3439), .Z(n2707) );
  CIVX2 U5431 ( .A(n2707), .Z(n2710) );
  CANR2X1 U5432 ( .A(n3435), .B(\m6.addrM64 [36]), .C(\m3.addrM64 [36]), .D(
        n3361), .Z(n2709) );
  CANR2X1 U5433 ( .A(n3436), .B(\m2.addrM64 [36]), .C(\m0.addrM64 [36]), .D(
        n3434), .Z(n2708) );
  CND4X2 U5434 ( .A(n2711), .B(n2710), .C(n2709), .D(n2708), .Z(n4124) );
  CAN2XL U5435 ( .A(\s6.addr [17]), .B(n4124), .Z(\s6.addr [36]) );
  CANR2X1 U5436 ( .A(n3431), .B(\m1.addrM64 [28]), .C(\m3.addrM64 [28]), .D(
        n3371), .Z(n2719) );
  CNR2IX1 U5437 ( .B(\m5.addrM64 [28]), .A(n3432), .Z(n2712) );
  CANR1X1 U5438 ( .A(n3434), .B(\m0.addrM64 [28]), .C(n2712), .Z(n2718) );
  CND2X1 U5439 ( .A(n3435), .B(\m6.addrM64 [28]), .Z(n2714) );
  CND2X1 U5440 ( .A(n3436), .B(\m2.addrM64 [28]), .Z(n2713) );
  CND2X1 U5441 ( .A(n2714), .B(n2713), .Z(n2716) );
  CNR2IX1 U5442 ( .B(\m4.addrM64 [28]), .A(n3439), .Z(n2715) );
  CNR2X1 U5443 ( .A(n2716), .B(n2715), .Z(n2717) );
  CND3X2 U5444 ( .A(n2719), .B(n2718), .C(n2717), .Z(n4133) );
  CAN2XL U5445 ( .A(\s6.addr [17]), .B(n4133), .Z(\s6.addr [28]) );
  CAN2XL U5446 ( .A(\s6.addr [17]), .B(n4128), .Z(\s6.addr [21]) );
  CNR2X4 U5447 ( .A(n2721), .B(n2720), .Z(n2722) );
  CIVX8 U5448 ( .A(n2722), .Z(n3453) );
  CIVX12 U5449 ( .A(n3453), .Z(\s1.en ) );
  CAOR2X1 U5450 ( .A(n4090), .B(\s1.dbus_out [39]), .C(n4094), .D(
        \s7.dbus_out [39]), .Z(n2742) );
  CIVX2 U5451 ( .A(n4335), .Z(n2723) );
  CND2X2 U5452 ( .A(n2724), .B(n2723), .Z(n2725) );
  CIVX2 U5453 ( .A(n2725), .Z(n2726) );
  CND2X2 U5454 ( .A(n2727), .B(n2726), .Z(n2739) );
  CIVX1 U5455 ( .A(n2729), .Z(n2730) );
  CND4X1 U5456 ( .A(n2731), .B(n2730), .C(n2762), .D(n3405), .Z(n2733) );
  CND3X4 U5457 ( .A(n2739), .B(n2738), .C(n2737), .Z(n3457) );
  CIVX8 U5458 ( .A(n2740), .Z(\s2.addr[16] ) );
  CAOR2XL U5459 ( .A(\c1.Breset ), .B(data_stm_d[39]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [39]), .Z(n2741) );
  CANR3XL U5460 ( .A(\s6.addr [17]), .B(\s6.dbus_out [39]), .C(n2742), .D(
        n2741), .Z(n2804) );
  CIVX8 U5461 ( .A(n3416), .Z(n4050) );
  CND2XL U5462 ( .A(n4098), .B(\s10.dbus_out [39]), .Z(n2749) );
  CNIVX1 U5463 ( .A(\s4.en ), .Z(n4077) );
  CANR2XL U5464 ( .A(n4078), .B(\s5.dbus_out [39]), .C(n4077), .D(
        \s4.dbus_out [39]), .Z(n2748) );
  CIVX16 U5465 ( .A(n3406), .Z(\s14.addr [11]) );
  CNIVX1 U5466 ( .A(\s14.addr [11]), .Z(n4100) );
  CNIVX2 U5467 ( .A(\s12.addr[11] ), .Z(n4099) );
  CANR2X1 U5468 ( .A(n4100), .B(\s14.dbus_out [39]), .C(\s12.dbus_out [39]), 
        .D(n4099), .Z(n2747) );
  CNR2X4 U5469 ( .A(n2744), .B(n2743), .Z(n2745) );
  CIVX8 U5470 ( .A(n2745), .Z(n3449) );
  CIVX16 U5471 ( .A(n3449), .Z(\s3.addr[9] ) );
  CND2XL U5472 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [39]), .Z(n2746) );
  CAN4X1 U5473 ( .A(n2749), .B(n2748), .C(n2747), .D(n2746), .Z(n2803) );
  CNIVX1 U5474 ( .A(\s11.addr[17] ), .Z(n4108) );
  CNR2X1 U5475 ( .A(n2750), .B(n2780), .Z(n2752) );
  CND2X1 U5476 ( .A(n2754), .B(n3485), .Z(n2757) );
  CIVX2 U5477 ( .A(n2755), .Z(n2756) );
  CND2X2 U5478 ( .A(n2759), .B(n2758), .Z(n2769) );
  CIVX2 U5479 ( .A(n2760), .Z(n2767) );
  CNR2X1 U5480 ( .A(n2761), .B(n3405), .Z(n2764) );
  CND3X2 U5481 ( .A(n2765), .B(n2764), .C(n2763), .Z(n2766) );
  CNR2X4 U5482 ( .A(n2767), .B(n2766), .Z(n2768) );
  CND2X4 U5483 ( .A(n2769), .B(n2768), .Z(n2770) );
  CIVX12 U5484 ( .A(n2770), .Z(n4188) );
  CAOR2XL U5485 ( .A(\s9.dbus_out [39]), .B(\s9.addr[8] ), .C(\s0.addr [14]), 
        .D(\s0.dbus_out [39]), .Z(n2771) );
  CANR1XL U5486 ( .A(n4108), .B(\s11.dbus_out [39]), .C(n2771), .Z(n2802) );
  CND3X1 U5487 ( .A(n3476), .B(n2772), .C(n4330), .Z(n2779) );
  CIVX1 U5488 ( .A(n2775), .Z(n2776) );
  COND1X2 U5489 ( .A(n2777), .B(n2776), .C(n3476), .Z(n2778) );
  CND3X2 U5490 ( .A(n1847), .B(n2784), .C(n2783), .Z(n2787) );
  CNR3X2 U5491 ( .A(n2787), .B(n2786), .C(n2785), .Z(n2799) );
  CND2X1 U5492 ( .A(n2794), .B(n2793), .Z(n2795) );
  CND3X2 U5493 ( .A(n2797), .B(n2796), .C(n2795), .Z(n2798) );
  CND3X4 U5494 ( .A(n2800), .B(n2799), .C(n2798), .Z(n3410) );
  CIVX16 U5495 ( .A(n2223), .Z(\s8.en ) );
  CANR2X1 U5496 ( .A(n4110), .B(\s13.dbus_out [39]), .C(n4085), .D(
        \s8.dbus_out [39]), .Z(n2801) );
  CND4XL U5497 ( .A(n2804), .B(n2803), .C(n2802), .D(n2801), .Z(n1715) );
  CAOR2X1 U5498 ( .A(n4095), .B(\s1.dbus_out [8]), .C(n4072), .D(
        \s7.dbus_out [8]), .Z(n2806) );
  CAOR2XL U5499 ( .A(\c1.Breset ), .B(data_stm_d[8]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [8]), .Z(n2805) );
  CANR3XL U5500 ( .A(\s6.addr [17]), .B(\s6.dbus_out [8]), .C(n2806), .D(n2805), .Z(n2821) );
  CANR1X4 U5501 ( .A(n2809), .B(n2808), .C(n2807), .Z(n2810) );
  CIVX8 U5502 ( .A(n2810), .Z(n3378) );
  CNR2IX1 U5503 ( .B(\s10.dbus_out [8]), .A(n4076), .Z(n2811) );
  CIVX2 U5504 ( .A(n2811), .Z(n2816) );
  CIVX4 U5505 ( .A(n2812), .Z(n5445) );
  CANR2XL U5506 ( .A(n4078), .B(\s5.dbus_out [8]), .C(n4077), .D(
        \s4.dbus_out [8]), .Z(n2815) );
  CANR2X1 U5507 ( .A(n4100), .B(\s14.dbus_out [8]), .C(\s12.dbus_out [8]), .D(
        n4099), .Z(n2814) );
  CND2XL U5508 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [8]), .Z(n2813) );
  CAN4X1 U5509 ( .A(n2816), .B(n2815), .C(n2814), .D(n2813), .Z(n2820) );
  CNIVX1 U5510 ( .A(\s11.en ), .Z(n4093) );
  CAOR2XL U5511 ( .A(\s9.dbus_out [8]), .B(\s9.addr[8] ), .C(\s0.en ), .D(
        \s0.dbus_out [8]), .Z(n2817) );
  CANR1XL U5512 ( .A(n4093), .B(\s11.dbus_out [8]), .C(n2817), .Z(n2819) );
  CANR2X1 U5513 ( .A(n4110), .B(\s13.dbus_out [8]), .C(n4109), .D(
        \s8.dbus_out [8]), .Z(n2818) );
  CND4XL U5514 ( .A(n2821), .B(n2820), .C(n2819), .D(n2818), .Z(n1746) );
  CAOR2XL U5515 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [0]), .C(n4072), .D(
        \s7.dbus_out [0]), .Z(n2823) );
  CAOR2XL U5516 ( .A(data_stm_d[0]), .B(\c1.Breset ), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [0]), .Z(n2822) );
  CANR3XL U5517 ( .A(n4062), .B(\s6.dbus_out [0]), .C(n2823), .D(n2822), .Z(
        n2832) );
  CND2X1 U5518 ( .A(n4098), .B(\s10.dbus_out [0]), .Z(n2827) );
  CANR2XL U5519 ( .A(n4078), .B(\s5.dbus_out [0]), .C(n4077), .D(
        \s4.dbus_out [0]), .Z(n2826) );
  CANR2XL U5520 ( .A(n4092), .B(\s14.dbus_out [0]), .C(\s12.dbus_out [0]), .D(
        \s12.addr[10] ), .Z(n2825) );
  CND2XL U5521 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [0]), .Z(n2824) );
  CAN4X1 U5522 ( .A(n2827), .B(n2826), .C(n2825), .D(n2824), .Z(n2831) );
  CIVX20 U5523 ( .A(n3298), .Z(\s9.addr[16] ) );
  CAOR2XL U5524 ( .A(\s9.dbus_out [0]), .B(\s9.addr[16] ), .C(n3940), .D(
        \s0.dbus_out [0]), .Z(n2828) );
  CANR1XL U5525 ( .A(n4108), .B(\s11.dbus_out [0]), .C(n2828), .Z(n2830) );
  CANR2XL U5526 ( .A(n4110), .B(\s13.dbus_out [0]), .C(n4085), .D(
        \s8.dbus_out [0]), .Z(n2829) );
  CND4XL U5527 ( .A(n2832), .B(n2831), .C(n2830), .D(n2829), .Z(n1754) );
  CNR2IX1 U5528 ( .B(\m5.addrM64 [46]), .A(n3432), .Z(n2833) );
  CNR2IX1 U5529 ( .B(\m4.addrM64 [46]), .A(n3439), .Z(n2834) );
  CIVX2 U5530 ( .A(n2834), .Z(n2838) );
  CANR2X1 U5531 ( .A(n3361), .B(\m3.addrM64 [46]), .C(\m6.addrM64 [46]), .D(
        n3435), .Z(n2837) );
  CAN2X1 U5532 ( .A(n3436), .B(\m2.addrM64 [46]), .Z(n2835) );
  CND4X2 U5533 ( .A(n2839), .B(n2838), .C(n2837), .D(n2836), .Z(n4136) );
  CAN2XL U5534 ( .A(\s6.addr [17]), .B(n4136), .Z(\s6.addr [46]) );
  CND2X1 U5535 ( .A(n3420), .B(\m3.addrM64 [44]), .Z(n2842) );
  CND2X1 U5536 ( .A(n3434), .B(\m0.addrM64 [44]), .Z(n2841) );
  CND2X1 U5537 ( .A(n3431), .B(\m1.addrM64 [44]), .Z(n2840) );
  CAN3X2 U5538 ( .A(n2842), .B(n2841), .C(n2840), .Z(n2850) );
  CIVX2 U5539 ( .A(\m5.addrM64 [44]), .Z(n2844) );
  CND2X1 U5540 ( .A(n3435), .B(\m6.addrM64 [44]), .Z(n2843) );
  CND2X1 U5541 ( .A(n3436), .B(\m2.addrM64 [44]), .Z(n2846) );
  CND2XL U5542 ( .A(n3424), .B(\m4.addrM64 [44]), .Z(n2845) );
  CND2X1 U5543 ( .A(n2846), .B(n2845), .Z(n2847) );
  CNR2X1 U5544 ( .A(n2848), .B(n2847), .Z(n2849) );
  CND2X2 U5545 ( .A(n2850), .B(n2849), .Z(n3470) );
  CAN2XL U5546 ( .A(\s6.addr [17]), .B(n3470), .Z(\s6.addr [44]) );
  CND2XL U5547 ( .A(n3431), .B(\m1.addrM64 [33]), .Z(n2852) );
  CND2XL U5548 ( .A(n3436), .B(\m2.addrM64 [33]), .Z(n2851) );
  CND2X1 U5549 ( .A(n2852), .B(n2851), .Z(n2854) );
  CNR2IX1 U5550 ( .B(\m4.addrM64 [33]), .A(n3439), .Z(n2853) );
  CNR2X1 U5551 ( .A(n2854), .B(n2853), .Z(n2859) );
  CANR2X1 U5552 ( .A(n2855), .B(\m3.addrM64 [33]), .C(\m6.addrM64 [33]), .D(
        n3435), .Z(n2858) );
  CNR2IX1 U5553 ( .B(\m5.addrM64 [33]), .A(n3432), .Z(n2856) );
  CANR1X1 U5554 ( .A(n3434), .B(\m0.addrM64 [33]), .C(n2856), .Z(n2857) );
  CND3X2 U5555 ( .A(n2859), .B(n2858), .C(n2857), .Z(n4179) );
  CAN2XL U5556 ( .A(\s6.addr [17]), .B(n4179), .Z(\s6.addr [33]) );
  CAN2XL U5557 ( .A(\s6.addr [17]), .B(n4134), .Z(\s6.addr [29]) );
  CNR2IX1 U5558 ( .B(\m4.addrM64 [26]), .A(n3439), .Z(n2860) );
  CNR2X1 U5559 ( .A(n2861), .B(n2860), .Z(n2866) );
  CANR2X1 U5560 ( .A(n3137), .B(\m3.addrM64 [26]), .C(\m6.addrM64 [26]), .D(
        n3435), .Z(n2865) );
  CND2X1 U5561 ( .A(n3434), .B(\m0.addrM64 [26]), .Z(n2863) );
  CNR2IX1 U5562 ( .B(\m5.addrM64 [26]), .A(n3432), .Z(n2862) );
  CNR2IX1 U5563 ( .B(n2863), .A(n2862), .Z(n2864) );
  CND3X2 U5564 ( .A(n2866), .B(n2865), .C(n2864), .Z(n4195) );
  CAN2XL U5565 ( .A(\s6.addr [17]), .B(n4195), .Z(\s6.addr [26]) );
  CND2X1 U5566 ( .A(n1842), .B(\m3.DoutM [27]), .Z(n2869) );
  CND2X1 U5567 ( .A(n3434), .B(\m0.DoutM [27]), .Z(n2868) );
  CND2X1 U5568 ( .A(n3431), .B(\m1.DoutM [27]), .Z(n2867) );
  CAN3X2 U5569 ( .A(n2869), .B(n2868), .C(n2867), .Z(n2875) );
  CIVX2 U5570 ( .A(\m5.DoutM [27]), .Z(n2871) );
  CND2X1 U5571 ( .A(n3435), .B(\m6.DoutM [27]), .Z(n2870) );
  CNR2X1 U5572 ( .A(n2873), .B(n2872), .Z(n2874) );
  CND2X2 U5573 ( .A(n2875), .B(n2874), .Z(n3460) );
  CAN2XL U5574 ( .A(\s6.addr [17]), .B(n3460), .Z(\s6.SbusIn [27]) );
  CND2X1 U5575 ( .A(n3434), .B(\m0.DoutM [29]), .Z(n2877) );
  CND2XL U5576 ( .A(n3436), .B(\m2.DoutM [29]), .Z(n2876) );
  CND2X1 U5577 ( .A(n2877), .B(n2876), .Z(n2881) );
  CIVX2 U5578 ( .A(\m5.DoutM [29]), .Z(n2879) );
  CND2X1 U5579 ( .A(n3435), .B(\m6.DoutM [29]), .Z(n2878) );
  CNR2X1 U5580 ( .A(n2881), .B(n2880), .Z(n2885) );
  CANR2X1 U5581 ( .A(n3431), .B(\m1.DoutM [29]), .C(\m3.DoutM [29]), .D(n3289), 
        .Z(n2884) );
  CNR2IX1 U5582 ( .B(\m4.DoutM [29]), .A(n3439), .Z(n2882) );
  CIVX2 U5583 ( .A(n2882), .Z(n2883) );
  CAN2XL U5584 ( .A(\s6.addr [17]), .B(n4197), .Z(\s6.SbusIn [29]) );
  CND2X1 U5585 ( .A(n3431), .B(\m1.DoutM [9]), .Z(n2887) );
  CND2XL U5586 ( .A(n3436), .B(\m2.DoutM [9]), .Z(n2886) );
  CND2X1 U5587 ( .A(n2887), .B(n2886), .Z(n2889) );
  CNR2IX1 U5588 ( .B(\m4.DoutM [9]), .A(n3439), .Z(n2888) );
  CNR2X1 U5589 ( .A(n2889), .B(n2888), .Z(n2893) );
  CANR2X1 U5590 ( .A(n3420), .B(\m3.DoutM [9]), .C(\m6.DoutM [9]), .D(n3435), 
        .Z(n2892) );
  CNR2IX1 U5591 ( .B(\m5.DoutM [9]), .A(n3432), .Z(n2890) );
  CANR1X1 U5592 ( .A(n3434), .B(\m0.DoutM [9]), .C(n2890), .Z(n2891) );
  CND3X2 U5593 ( .A(n2893), .B(n2892), .C(n2891), .Z(n4193) );
  CAN2XL U5594 ( .A(\s6.addr [17]), .B(n4193), .Z(\s6.SbusIn [9]) );
  CIVX1 U5595 ( .A(\c1.Breset ), .Z(n5518) );
  CAOR2XL U5596 ( .A(n4090), .B(\s1.dbus_out [14]), .C(n4094), .D(
        \s7.dbus_out [14]), .Z(n2895) );
  CAOR2XL U5597 ( .A(\c1.Breset ), .B(data_stm_d[14]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [14]), .Z(n2894) );
  CANR3XL U5598 ( .A(n4062), .B(\s6.dbus_out [14]), .C(n2895), .D(n2894), .Z(
        n2904) );
  CND2X1 U5599 ( .A(n4098), .B(\s10.dbus_out [14]), .Z(n2899) );
  CNIVX1 U5600 ( .A(\s4.addr[14] ), .Z(n4091) );
  CANR2XL U5601 ( .A(n4078), .B(\s5.dbus_out [14]), .C(n4091), .D(
        \s4.dbus_out [14]), .Z(n2898) );
  CANR2X1 U5602 ( .A(n4092), .B(\s14.dbus_out [14]), .C(\s12.dbus_out [14]), 
        .D(n4099), .Z(n2897) );
  CND2X1 U5603 ( .A(n4101), .B(\s3.dbus_out [14]), .Z(n2896) );
  CAN4X1 U5604 ( .A(n2899), .B(n2898), .C(n2897), .D(n2896), .Z(n2903) );
  CIVX16 U5605 ( .A(n3298), .Z(\s9.addr[7] ) );
  CAOR2XL U5606 ( .A(\s9.dbus_out [14]), .B(n5590), .C(n4083), .D(
        \s0.dbus_out [14]), .Z(n2900) );
  CANR1XL U5607 ( .A(n4093), .B(\s11.dbus_out [14]), .C(n2900), .Z(n2902) );
  CANR2X1 U5608 ( .A(n4110), .B(\s13.dbus_out [14]), .C(n4085), .D(
        \s8.dbus_out [14]), .Z(n2901) );
  CND4XL U5609 ( .A(n2904), .B(n2903), .C(n2902), .D(n2901), .Z(n1740) );
  CND2X1 U5610 ( .A(n3420), .B(\m3.addrM64 [34]), .Z(n2907) );
  CND2XL U5611 ( .A(n3434), .B(\m0.addrM64 [34]), .Z(n2906) );
  CND2X1 U5612 ( .A(n3431), .B(\m1.addrM64 [34]), .Z(n2905) );
  CAN3X2 U5613 ( .A(n2907), .B(n2906), .C(n2905), .Z(n2915) );
  CIVX2 U5614 ( .A(\m5.addrM64 [34]), .Z(n2909) );
  CND2X1 U5615 ( .A(n3435), .B(\m6.addrM64 [34]), .Z(n2908) );
  CIVX2 U5616 ( .A(\m4.addrM64 [34]), .Z(n2911) );
  CND2X1 U5617 ( .A(n3436), .B(\m2.addrM64 [34]), .Z(n2910) );
  CNR2X1 U5618 ( .A(n2913), .B(n2912), .Z(n2914) );
  CND2X2 U5619 ( .A(n2915), .B(n2914), .Z(n4131) );
  CAN2XL U5620 ( .A(n1844), .B(n4131), .Z(\s5.addr [34]) );
  CND2XL U5621 ( .A(n3431), .B(\m1.addrM64 [31]), .Z(n2917) );
  CND2XL U5622 ( .A(n3436), .B(\m2.addrM64 [31]), .Z(n2916) );
  CND2X1 U5623 ( .A(n2917), .B(n2916), .Z(n2919) );
  CNR2IX1 U5624 ( .B(\m4.addrM64 [31]), .A(n3439), .Z(n2918) );
  CNR2X1 U5625 ( .A(n2919), .B(n2918), .Z(n2923) );
  CANR2X1 U5626 ( .A(n3361), .B(\m3.addrM64 [31]), .C(\m6.addrM64 [31]), .D(
        n3435), .Z(n2922) );
  CNR2IX1 U5627 ( .B(\m5.addrM64 [31]), .A(n3432), .Z(n2920) );
  CANR1X1 U5628 ( .A(n3434), .B(\m0.addrM64 [31]), .C(n2920), .Z(n2921) );
  CND3X2 U5629 ( .A(n2923), .B(n2922), .C(n2921), .Z(n4160) );
  CAN2XL U5630 ( .A(n5445), .B(n4160), .Z(\s5.addr [31]) );
  CANR2X1 U5631 ( .A(n3431), .B(\m1.addrM64 [51]), .C(\m3.addrM64 [51]), .D(
        n3090), .Z(n2931) );
  CNR2IX1 U5632 ( .B(\m5.addrM64 [51]), .A(n3432), .Z(n2924) );
  CANR1X1 U5633 ( .A(n3434), .B(\m0.addrM64 [51]), .C(n2924), .Z(n2930) );
  CND2X1 U5634 ( .A(n3435), .B(\m6.addrM64 [51]), .Z(n2926) );
  CND2X1 U5635 ( .A(n3436), .B(\m2.addrM64 [51]), .Z(n2925) );
  CND2X1 U5636 ( .A(n2926), .B(n2925), .Z(n2928) );
  CNR2IX1 U5637 ( .B(\m4.addrM64 [51]), .A(n3439), .Z(n2927) );
  CNR2X1 U5638 ( .A(n2928), .B(n2927), .Z(n2929) );
  CND3X2 U5639 ( .A(n2931), .B(n2930), .C(n2929), .Z(n4165) );
  CAN2XL U5640 ( .A(n4405), .B(n4165), .Z(\s5.addr [51]) );
  CND2X1 U5641 ( .A(n3431), .B(\m1.addrM64 [27]), .Z(n2933) );
  CND2XL U5642 ( .A(n3436), .B(\m2.addrM64 [27]), .Z(n2932) );
  CND2X1 U5643 ( .A(n2933), .B(n2932), .Z(n2935) );
  CNR2IX1 U5644 ( .B(\m4.addrM64 [27]), .A(n3439), .Z(n2934) );
  CNR2X1 U5645 ( .A(n2935), .B(n2934), .Z(n2939) );
  CANR2X1 U5646 ( .A(n3090), .B(\m3.addrM64 [27]), .C(\m6.addrM64 [27]), .D(
        n3435), .Z(n2938) );
  CNR2IX1 U5647 ( .B(\m5.addrM64 [27]), .A(n3432), .Z(n2936) );
  CANR1X1 U5648 ( .A(n3434), .B(\m0.addrM64 [27]), .C(n2936), .Z(n2937) );
  CND3X2 U5649 ( .A(n2939), .B(n2938), .C(n2937), .Z(n3467) );
  CAN2XL U5650 ( .A(n4405), .B(n3467), .Z(\s5.addr [27]) );
  CANR2X1 U5651 ( .A(n3431), .B(\m1.addrM64 [59]), .C(\m3.addrM64 [59]), .D(
        n3361), .Z(n2946) );
  CND2X1 U5652 ( .A(n3434), .B(\m0.addrM64 [59]), .Z(n2941) );
  CNR2IX1 U5653 ( .B(\m5.addrM64 [59]), .A(n3432), .Z(n2940) );
  CNR2IX1 U5654 ( .B(n2941), .A(n2940), .Z(n2945) );
  CAN2XL U5655 ( .A(n3424), .B(\m4.addrM64 [59]), .Z(n2942) );
  CNR2X1 U5656 ( .A(n2943), .B(n2942), .Z(n2944) );
  CAN2XL U5657 ( .A(n4405), .B(n3477), .Z(\s5.addr [59]) );
  CNR2IX1 U5658 ( .B(\m5.addrM64 [62]), .A(n3432), .Z(n2947) );
  CND2X1 U5659 ( .A(n3424), .B(\m4.addrM64 [62]), .Z(n2950) );
  CANR2X1 U5660 ( .A(n3137), .B(\m3.addrM64 [62]), .C(\m6.addrM64 [62]), .D(
        n3435), .Z(n2949) );
  CANR2X1 U5661 ( .A(n3436), .B(\m2.addrM64 [62]), .C(\m0.addrM64 [62]), .D(
        n3434), .Z(n2948) );
  CND4X2 U5662 ( .A(n2951), .B(n2950), .C(n2949), .D(n2948), .Z(n3479) );
  CAN2XL U5663 ( .A(n1844), .B(n3479), .Z(\s5.addr [62]) );
  CAN2XL U5664 ( .A(n5445), .B(n3483), .Z(\s5.SbusIn [23]) );
  CAN2XL U5665 ( .A(n4405), .B(n3465), .Z(\s5.SbusIn [11]) );
  CANR2X1 U5666 ( .A(n3431), .B(\m1.DoutM [24]), .C(\m3.DoutM [24]), .D(n3420), 
        .Z(n2959) );
  CNR2IX1 U5667 ( .B(\m5.DoutM [24]), .A(n3432), .Z(n2952) );
  CND2X1 U5668 ( .A(n3435), .B(\m6.DoutM [24]), .Z(n2954) );
  CND2X1 U5669 ( .A(n3436), .B(\m2.DoutM [24]), .Z(n2953) );
  CND2X1 U5670 ( .A(n2954), .B(n2953), .Z(n2956) );
  CNR2IX1 U5671 ( .B(\m4.DoutM [24]), .A(n3439), .Z(n2955) );
  CNR2X1 U5672 ( .A(n2956), .B(n2955), .Z(n2957) );
  CND3X2 U5673 ( .A(n2959), .B(n2958), .C(n2957), .Z(n4149) );
  CAN2XL U5674 ( .A(\s6.addr [17]), .B(n4149), .Z(\s6.SbusIn [24]) );
  CND2X1 U5675 ( .A(n3434), .B(\m0.addrM64 [49]), .Z(n2961) );
  CND2XL U5676 ( .A(n3436), .B(\m2.addrM64 [49]), .Z(n2960) );
  CND2X1 U5677 ( .A(n2961), .B(n2960), .Z(n2965) );
  CIVX2 U5678 ( .A(\m5.addrM64 [49]), .Z(n2963) );
  CND2X1 U5679 ( .A(n3435), .B(\m6.addrM64 [49]), .Z(n2962) );
  CNR2X1 U5680 ( .A(n2965), .B(n2964), .Z(n2969) );
  CANR2X1 U5681 ( .A(n3431), .B(\m1.addrM64 [49]), .C(\m3.addrM64 [49]), .D(
        n3420), .Z(n2968) );
  CNR2IX1 U5682 ( .B(\m4.addrM64 [49]), .A(n3439), .Z(n2966) );
  CIVX2 U5683 ( .A(n2966), .Z(n2967) );
  CAN2XL U5684 ( .A(\s6.addr [17]), .B(n4155), .Z(\s6.addr [49]) );
  CANR2X1 U5685 ( .A(n3431), .B(\m1.addrM64 [54]), .C(\m3.addrM64 [54]), .D(
        n3361), .Z(n2977) );
  CNR2IX1 U5686 ( .B(\m5.addrM64 [54]), .A(n3432), .Z(n2970) );
  CANR1X1 U5687 ( .A(n3434), .B(\m0.addrM64 [54]), .C(n2970), .Z(n2976) );
  CND2X1 U5688 ( .A(n3435), .B(\m6.addrM64 [54]), .Z(n2972) );
  CND2X1 U5689 ( .A(n3436), .B(\m2.addrM64 [54]), .Z(n2971) );
  CND2X1 U5690 ( .A(n2972), .B(n2971), .Z(n2974) );
  CAN2XL U5691 ( .A(n3424), .B(\m4.addrM64 [54]), .Z(n2973) );
  CNR2X1 U5692 ( .A(n2974), .B(n2973), .Z(n2975) );
  CND3X2 U5693 ( .A(n2977), .B(n2976), .C(n2975), .Z(n4148) );
  CAN2XL U5694 ( .A(\s6.addr [17]), .B(n4148), .Z(\s6.addr [54]) );
  CIVX8 U5695 ( .A(\m4.ack ), .Z(n2978) );
  CNR2XL U5696 ( .A(n2978), .B(n5564), .Z(\m4.MinData [41]) );
  CNR2XL U5697 ( .A(n2978), .B(n5563), .Z(\m4.MinData [40]) );
  CNR2XL U5698 ( .A(n2978), .B(n5562), .Z(\m4.MinData [39]) );
  CNR2XL U5699 ( .A(n2978), .B(n5561), .Z(\m4.MinData [38]) );
  CNR2XL U5700 ( .A(n2978), .B(n5560), .Z(\m4.MinData [37]) );
  CNR2XL U5701 ( .A(n2978), .B(n5559), .Z(\m4.MinData [36]) );
  CNR2XL U5702 ( .A(n2978), .B(n5558), .Z(\m4.MinData [35]) );
  CNR2XL U5703 ( .A(n2978), .B(n5557), .Z(\m4.MinData [34]) );
  CNR2XL U5704 ( .A(n2978), .B(n5556), .Z(\m4.MinData [33]) );
  CNR2XL U5705 ( .A(n2978), .B(n5555), .Z(\m4.MinData [32]) );
  CNR2XL U5706 ( .A(n2978), .B(n5554), .Z(\m4.MinData [31]) );
  CNR2XL U5707 ( .A(n2978), .B(n5553), .Z(\m4.MinData [30]) );
  CNR2XL U5708 ( .A(n2978), .B(n5552), .Z(\m4.MinData [29]) );
  CNR2XL U5709 ( .A(n2978), .B(n5551), .Z(\m4.MinData [28]) );
  CNR2XL U5710 ( .A(n2978), .B(n5565), .Z(\m4.MinData [42]) );
  CNR2XL U5711 ( .A(n2978), .B(n5566), .Z(\m4.MinData [43]) );
  CNR2XL U5712 ( .A(n2978), .B(n5567), .Z(\m4.MinData [44]) );
  CNR2XL U5713 ( .A(n2978), .B(n5568), .Z(\m4.MinData [45]) );
  CNR2XL U5714 ( .A(n2978), .B(n5569), .Z(\m4.MinData [46]) );
  CNR2XL U5715 ( .A(n2978), .B(n5570), .Z(\m4.MinData [47]) );
  CNR2XL U5716 ( .A(n2978), .B(n5571), .Z(\m4.MinData [48]) );
  CNR2XL U5717 ( .A(n2978), .B(n5572), .Z(\m4.MinData [49]) );
  CNR2XL U5718 ( .A(n2978), .B(n5574), .Z(\m4.MinData [50]) );
  CNR2XL U5719 ( .A(n2978), .B(n5575), .Z(\m4.MinData [51]) );
  CNR2XL U5720 ( .A(n2978), .B(n5576), .Z(\m4.MinData [52]) );
  CNR2XL U5721 ( .A(n2978), .B(n5577), .Z(\m4.MinData [53]) );
  CNR2XL U5722 ( .A(n2978), .B(n5578), .Z(\m4.MinData [54]) );
  CNR2XL U5723 ( .A(n2978), .B(n5579), .Z(\m4.MinData [55]) );
  CNR2XL U5724 ( .A(n2978), .B(n5580), .Z(\m4.MinData [56]) );
  CNR2XL U5725 ( .A(n2978), .B(n5581), .Z(\m4.MinData [57]) );
  CNR2XL U5726 ( .A(n2978), .B(n5587), .Z(\m4.MinData [63]) );
  CNR2XL U5727 ( .A(n2978), .B(n5582), .Z(\m4.MinData [58]) );
  CNR2XL U5728 ( .A(n2978), .B(n5583), .Z(\m4.MinData [59]) );
  CNR2XL U5729 ( .A(n2978), .B(n5584), .Z(\m4.MinData [60]) );
  CNR2XL U5730 ( .A(n2978), .B(n5586), .Z(\m4.MinData [62]) );
  CNR2XL U5731 ( .A(n2978), .B(n5585), .Z(\m4.MinData [61]) );
  CNR2XL U5732 ( .A(n2978), .B(n5539), .Z(\m4.MinData [16]) );
  CNR2XL U5733 ( .A(n2978), .B(n5528), .Z(\m4.MinData [5]) );
  CNR2XL U5734 ( .A(n2978), .B(n5550), .Z(\m4.MinData [27]) );
  CNR2XL U5735 ( .A(n2978), .B(n5538), .Z(\m4.MinData [15]) );
  CNR2XL U5736 ( .A(n2978), .B(n5540), .Z(\m4.MinData [17]) );
  CNR2XL U5737 ( .A(n2978), .B(n5549), .Z(\m4.MinData [26]) );
  CNR2XL U5738 ( .A(n2978), .B(n5523), .Z(\m4.MinData [0]) );
  CNR2XL U5739 ( .A(n2978), .B(n5524), .Z(\m4.MinData [1]) );
  CNR2XL U5740 ( .A(n2978), .B(n5548), .Z(\m4.MinData [25]) );
  CNR2XL U5741 ( .A(n2978), .B(n5525), .Z(\m4.MinData [2]) );
  CNR2XL U5742 ( .A(n2978), .B(n5526), .Z(\m4.MinData [3]) );
  CNR2XL U5743 ( .A(n2978), .B(n5532), .Z(\m4.MinData [9]) );
  CNR2XL U5744 ( .A(n2978), .B(n5547), .Z(\m4.MinData [24]) );
  CNR2XL U5745 ( .A(n2978), .B(n5527), .Z(\m4.MinData [4]) );
  CNR2XL U5746 ( .A(n2978), .B(n5533), .Z(\m4.MinData [10]) );
  CNR2XL U5747 ( .A(n2978), .B(n5546), .Z(\m4.MinData [23]) );
  CNR2XL U5748 ( .A(n2978), .B(n5534), .Z(\m4.MinData [11]) );
  CNR2XL U5749 ( .A(n2978), .B(n5537), .Z(\m4.MinData [14]) );
  CNR2XL U5750 ( .A(n2978), .B(n5529), .Z(\m4.MinData [6]) );
  CNR2XL U5751 ( .A(n2978), .B(n5536), .Z(\m4.MinData [13]) );
  CNR2XL U5752 ( .A(n2978), .B(n5541), .Z(\m4.MinData [18]) );
  CNR2XL U5753 ( .A(n2978), .B(n5530), .Z(\m4.MinData [7]) );
  CNR2XL U5754 ( .A(n2978), .B(n5545), .Z(\m4.MinData [22]) );
  CNR2XL U5755 ( .A(n2978), .B(n5535), .Z(\m4.MinData [12]) );
  CNR2XL U5756 ( .A(n2978), .B(n5531), .Z(\m4.MinData [8]) );
  CNR2XL U5757 ( .A(n2978), .B(n5544), .Z(\m4.MinData [21]) );
  CNR2XL U5758 ( .A(n2978), .B(n5542), .Z(\m4.MinData [19]) );
  CNR2XL U5759 ( .A(n2978), .B(n5543), .Z(\m4.MinData [20]) );
  CNR2XL U5760 ( .A(n2979), .B(n5530), .Z(\m5.MinData [7]) );
  CNR2XL U5761 ( .A(n2979), .B(n5542), .Z(\m5.MinData [19]) );
  CNR2XL U5762 ( .A(n2979), .B(n5569), .Z(\m5.MinData [46]) );
  CNR2XL U5763 ( .A(n2979), .B(n5568), .Z(\m5.MinData [45]) );
  CNR2XL U5764 ( .A(n2979), .B(n5566), .Z(\m5.MinData [43]) );
  CNR2XL U5765 ( .A(n2979), .B(n5539), .Z(\m5.MinData [16]) );
  CNR2XL U5766 ( .A(n2979), .B(n5531), .Z(\m5.MinData [8]) );
  CNR2XL U5767 ( .A(n2979), .B(n5540), .Z(\m5.MinData [17]) );
  CNR2XL U5768 ( .A(n2979), .B(n5564), .Z(\m5.MinData [41]) );
  CNR2XL U5769 ( .A(n2979), .B(n5565), .Z(\m5.MinData [42]) );
  CNR2XL U5770 ( .A(n2979), .B(n5567), .Z(\m5.MinData [44]) );
  CNR2XL U5771 ( .A(n2979), .B(n5541), .Z(\m5.MinData [18]) );
  CNR2XL U5772 ( .A(n2979), .B(n5576), .Z(\m5.MinData [52]) );
  CNR2XL U5773 ( .A(n2979), .B(n5528), .Z(\m5.MinData [5]) );
  CNR2XL U5774 ( .A(n2979), .B(n5577), .Z(\m5.MinData [53]) );
  CNR2XL U5775 ( .A(n2979), .B(n5562), .Z(\m5.MinData [39]) );
  CNR2XL U5776 ( .A(n2979), .B(n5534), .Z(\m5.MinData [11]) );
  CNR2XL U5777 ( .A(n2979), .B(n5575), .Z(\m5.MinData [51]) );
  CNR2XL U5778 ( .A(n2979), .B(n5527), .Z(\m5.MinData [4]) );
  CNR2XL U5779 ( .A(n2979), .B(n5578), .Z(\m5.MinData [54]) );
  CNR2XL U5780 ( .A(n2979), .B(n5563), .Z(\m5.MinData [40]) );
  CNR2XL U5781 ( .A(n2979), .B(n5574), .Z(\m5.MinData [50]) );
  CNR2XL U5782 ( .A(n2979), .B(n5579), .Z(\m5.MinData [55]) );
  CNR2XL U5783 ( .A(n2979), .B(n5580), .Z(\m5.MinData [56]) );
  CNR2XL U5784 ( .A(n2979), .B(n5529), .Z(\m5.MinData [6]) );
  CNR2XL U5785 ( .A(n2979), .B(n5535), .Z(\m5.MinData [12]) );
  CNR2XL U5786 ( .A(n2979), .B(n5581), .Z(\m5.MinData [57]) );
  CNR2XL U5787 ( .A(n2979), .B(n5582), .Z(\m5.MinData [58]) );
  CNR2XL U5788 ( .A(n2979), .B(n5526), .Z(\m5.MinData [3]) );
  CNR2XL U5789 ( .A(n2979), .B(n5583), .Z(\m5.MinData [59]) );
  CNR2XL U5790 ( .A(n2979), .B(n5584), .Z(\m5.MinData [60]) );
  CNR2XL U5791 ( .A(n2979), .B(n5572), .Z(\m5.MinData [49]) );
  CNR2XL U5792 ( .A(n2979), .B(n5585), .Z(\m5.MinData [61]) );
  CNR2XL U5793 ( .A(n2979), .B(n5586), .Z(\m5.MinData [62]) );
  CNR2XL U5794 ( .A(n2979), .B(n5536), .Z(\m5.MinData [13]) );
  CNR2XL U5795 ( .A(n2979), .B(n5525), .Z(\m5.MinData [2]) );
  CNR2XL U5796 ( .A(n2979), .B(n5587), .Z(\m5.MinData [63]) );
  CNR2XL U5797 ( .A(n2979), .B(n5524), .Z(\m5.MinData [1]) );
  CNR2XL U5798 ( .A(n2979), .B(n5533), .Z(\m5.MinData [10]) );
  CNR2XL U5799 ( .A(n2979), .B(n5523), .Z(\m5.MinData [0]) );
  CNR2XL U5800 ( .A(n2979), .B(n5571), .Z(\m5.MinData [48]) );
  CNR2XL U5801 ( .A(n2979), .B(n5537), .Z(\m5.MinData [14]) );
  CNR2XL U5802 ( .A(n2979), .B(n5538), .Z(\m5.MinData [15]) );
  CNR2XL U5803 ( .A(n2979), .B(n5570), .Z(\m5.MinData [47]) );
  CNR2XL U5804 ( .A(n2979), .B(n5561), .Z(\m5.MinData [38]) );
  CNR2XL U5805 ( .A(n2979), .B(n5532), .Z(\m5.MinData [9]) );
  CNR2XL U5806 ( .A(n2979), .B(n5546), .Z(\m5.MinData [23]) );
  CNR2XL U5807 ( .A(n2979), .B(n5551), .Z(\m5.MinData [28]) );
  CNR2XL U5808 ( .A(n2979), .B(n5557), .Z(\m5.MinData [34]) );
  CNR2XL U5809 ( .A(n2979), .B(n5559), .Z(\m5.MinData [36]) );
  CNR2XL U5810 ( .A(n2979), .B(n5547), .Z(\m5.MinData [24]) );
  CNR2XL U5811 ( .A(n2979), .B(n5558), .Z(\m5.MinData [35]) );
  CNR2XL U5812 ( .A(n2979), .B(n5548), .Z(\m5.MinData [25]) );
  CNR2XL U5813 ( .A(n2979), .B(n5549), .Z(\m5.MinData [26]) );
  CNR2XL U5814 ( .A(n2979), .B(n5550), .Z(\m5.MinData [27]) );
  CNR2XL U5815 ( .A(n2979), .B(n5554), .Z(\m5.MinData [31]) );
  CNR2XL U5816 ( .A(n2979), .B(n5560), .Z(\m5.MinData [37]) );
  CNR2XL U5817 ( .A(n2979), .B(n5543), .Z(\m5.MinData [20]) );
  CNR2XL U5818 ( .A(n2979), .B(n5553), .Z(\m5.MinData [30]) );
  CNR2XL U5819 ( .A(n2979), .B(n5544), .Z(\m5.MinData [21]) );
  CNR2XL U5820 ( .A(n2979), .B(n5555), .Z(\m5.MinData [32]) );
  CNR2XL U5821 ( .A(n2979), .B(n5556), .Z(\m5.MinData [33]) );
  CNR2XL U5822 ( .A(n2979), .B(n5552), .Z(\m5.MinData [29]) );
  CNR2XL U5823 ( .A(n2979), .B(n5545), .Z(\m5.MinData [22]) );
  CNR2XL U5824 ( .A(n3383), .B(n5538), .Z(\m1.MinData [15]) );
  CNR2XL U5825 ( .A(n3383), .B(n5536), .Z(\m1.MinData [13]) );
  CNR2XL U5826 ( .A(n3383), .B(n5537), .Z(\m1.MinData [14]) );
  CNR2XL U5827 ( .A(n3383), .B(n5534), .Z(\m1.MinData [11]) );
  CNR2XL U5828 ( .A(n3383), .B(n5539), .Z(\m1.MinData [16]) );
  CNR2XL U5829 ( .A(n3383), .B(n5531), .Z(\m1.MinData [8]) );
  CNR2XL U5830 ( .A(n3383), .B(n5540), .Z(\m1.MinData [17]) );
  CNR2XL U5831 ( .A(n3383), .B(n5529), .Z(\m1.MinData [6]) );
  CNR2XL U5832 ( .A(n3383), .B(n5532), .Z(\m1.MinData [9]) );
  CNR2XL U5833 ( .A(n3383), .B(n5541), .Z(\m1.MinData [18]) );
  CNR2XL U5834 ( .A(n3383), .B(n5535), .Z(\m1.MinData [12]) );
  CNR2XL U5835 ( .A(n3383), .B(n5533), .Z(\m1.MinData [10]) );
  CNR2XL U5836 ( .A(n3383), .B(n5542), .Z(\m1.MinData [19]) );
  CNR2XL U5837 ( .A(n3383), .B(n5543), .Z(\m1.MinData [20]) );
  CNR2XL U5838 ( .A(n3383), .B(n5544), .Z(\m1.MinData [21]) );
  CNR2XL U5839 ( .A(n3383), .B(n5528), .Z(\m1.MinData [5]) );
  CNR2XL U5840 ( .A(n3383), .B(n5546), .Z(\m1.MinData [23]) );
  CNR2XL U5841 ( .A(n3383), .B(n5547), .Z(\m1.MinData [24]) );
  CNR2XL U5842 ( .A(n3383), .B(n5549), .Z(\m1.MinData [26]) );
  CNR2XL U5843 ( .A(n3383), .B(n5550), .Z(\m1.MinData [27]) );
  CNR2XL U5844 ( .A(n3383), .B(n5552), .Z(\m1.MinData [29]) );
  CNR2XL U5845 ( .A(n3383), .B(n5553), .Z(\m1.MinData [30]) );
  CNR2XL U5846 ( .A(n3383), .B(n5555), .Z(\m1.MinData [32]) );
  CNR2XL U5847 ( .A(n3383), .B(n5556), .Z(\m1.MinData [33]) );
  CNR2XL U5848 ( .A(n3383), .B(n5558), .Z(\m1.MinData [35]) );
  CNR2XL U5849 ( .A(n3383), .B(n5560), .Z(\m1.MinData [37]) );
  CNR2XL U5850 ( .A(n3383), .B(n5561), .Z(\m1.MinData [38]) );
  CNR2XL U5851 ( .A(n3383), .B(n5586), .Z(\m1.MinData [62]) );
  CNR2XL U5852 ( .A(n3383), .B(n5585), .Z(\m1.MinData [61]) );
  CNR2XL U5853 ( .A(n3383), .B(n5564), .Z(\m1.MinData [41]) );
  CNR2XL U5854 ( .A(n3383), .B(n5565), .Z(\m1.MinData [42]) );
  CNR2XL U5855 ( .A(n3383), .B(n5583), .Z(\m1.MinData [59]) );
  CNR2XL U5856 ( .A(n3383), .B(n5567), .Z(\m1.MinData [44]) );
  CNR2XL U5857 ( .A(n3383), .B(n5568), .Z(\m1.MinData [45]) );
  CNR2XL U5858 ( .A(n3383), .B(n5581), .Z(\m1.MinData [57]) );
  CNR2XL U5859 ( .A(n3383), .B(n5571), .Z(\m1.MinData [48]) );
  CNR2XL U5860 ( .A(n3383), .B(n5580), .Z(\m1.MinData [56]) );
  CNR2XL U5861 ( .A(n3383), .B(n5572), .Z(\m1.MinData [49]) );
  CNR2XL U5862 ( .A(n3383), .B(n5574), .Z(\m1.MinData [50]) );
  CNR2XL U5863 ( .A(n3383), .B(n5576), .Z(\m1.MinData [52]) );
  CNR2XL U5864 ( .A(n3383), .B(n5577), .Z(\m1.MinData [53]) );
  CND2X4 U5865 ( .A(n3420), .B(n5518), .Z(n3379) );
  CIVX2 U5866 ( .A(n3379), .Z(\m3.ack ) );
  CNR2XL U5867 ( .A(n3383), .B(n5569), .Z(\m1.MinData [46]) );
  CNIVX4 U5868 ( .A(n3463), .Z(\s9.addr [15]) );
  CAN2X1 U5869 ( .A(\s7.en ), .B(n3478), .Z(\s7.addr [6]) );
  CNIVX4 U5870 ( .A(\s14.addr [11]), .Z(\s14.addr[16] ) );
  CAN2XL U5871 ( .A(n4405), .B(n4150), .Z(\s5.SbusIn [20]) );
  CAN2XL U5872 ( .A(n4405), .B(n3472), .Z(\s5.SbusIn [46]) );
  CAN2XL U5873 ( .A(n1844), .B(n4149), .Z(\s5.SbusIn [24]) );
  CAN2XL U5874 ( .A(n5445), .B(n4197), .Z(\s5.SbusIn [29]) );
  CAN2XL U5875 ( .A(\s6.addr [17]), .B(n4138), .Z(\s6.SbusIn [44]) );
  CAN2XL U5876 ( .A(\s6.addr [17]), .B(n4117), .Z(\s6.SbusIn [28]) );
  CAN2XL U5877 ( .A(\s6.addr [17]), .B(n4171), .Z(\s6.SbusIn [32]) );
  CNR2IX1 U5878 ( .B(\m5.DoutM [21]), .A(n3432), .Z(n2980) );
  CNR2IX1 U5879 ( .B(\m4.DoutM [21]), .A(n3439), .Z(n2981) );
  CIVX2 U5880 ( .A(n2981), .Z(n2984) );
  CANR2X1 U5881 ( .A(n3361), .B(\m3.DoutM [21]), .C(\m6.DoutM [21]), .D(n3435), 
        .Z(n2983) );
  CANR2X1 U5882 ( .A(n3434), .B(\m0.DoutM [21]), .C(n3436), .D(\m2.DoutM [21]), 
        .Z(n2982) );
  CND4X2 U5883 ( .A(n2985), .B(n2984), .C(n2983), .D(n2982), .Z(n4158) );
  CAN2XL U5884 ( .A(\s6.addr [17]), .B(n4158), .Z(\s6.SbusIn [21]) );
  CAN2XL U5885 ( .A(\s6.addr [17]), .B(n4237), .Z(\s6.SbusIn [35]) );
  CNR2IX1 U5886 ( .B(\m4.DoutM [36]), .A(n3439), .Z(n2986) );
  CNR2X1 U5887 ( .A(n2987), .B(n2986), .Z(n2991) );
  CANR2X1 U5888 ( .A(n3420), .B(\m3.DoutM [36]), .C(\m6.DoutM [36]), .D(n3435), 
        .Z(n2990) );
  CNR2IX1 U5889 ( .B(\m5.DoutM [36]), .A(n3432), .Z(n2988) );
  CND3X2 U5890 ( .A(n2991), .B(n2990), .C(n2989), .Z(n4215) );
  CAN2XL U5891 ( .A(\s6.addr [17]), .B(n4215), .Z(\s6.SbusIn [36]) );
  CAN2XL U5892 ( .A(\s6.addr [17]), .B(n4135), .Z(\s6.SbusIn [39]) );
  CNR2IX1 U5893 ( .B(\m4.DoutM [15]), .A(n3439), .Z(n2992) );
  CNR2X1 U5894 ( .A(n2993), .B(n2992), .Z(n2998) );
  CANR2X1 U5895 ( .A(n3289), .B(\m3.DoutM [15]), .C(\m6.DoutM [15]), .D(n3435), 
        .Z(n2997) );
  CND2X1 U5896 ( .A(n3434), .B(\m0.DoutM [15]), .Z(n2995) );
  CNR2IX1 U5897 ( .B(\m5.DoutM [15]), .A(n3432), .Z(n2994) );
  CNR2IX1 U5898 ( .B(n2995), .A(n2994), .Z(n2996) );
  CND3X2 U5899 ( .A(n2998), .B(n2997), .C(n2996), .Z(n4169) );
  CAN2XL U5900 ( .A(\s6.addr [17]), .B(n4169), .Z(\s6.SbusIn [15]) );
  CAN2XL U5901 ( .A(\s6.addr [17]), .B(n3467), .Z(\s6.addr [27]) );
  CND2X1 U5902 ( .A(n3431), .B(\m1.addrM64 [35]), .Z(n3000) );
  CND2XL U5903 ( .A(n3436), .B(\m2.addrM64 [35]), .Z(n2999) );
  CND2X1 U5904 ( .A(n3000), .B(n2999), .Z(n3002) );
  CNR2IX1 U5905 ( .B(\m4.addrM64 [35]), .A(n3439), .Z(n3001) );
  CNR2X1 U5906 ( .A(n3002), .B(n3001), .Z(n3006) );
  CANR2X1 U5907 ( .A(n3435), .B(\m6.addrM64 [35]), .C(\m3.addrM64 [35]), .D(
        n3420), .Z(n3005) );
  CNR2IX1 U5908 ( .B(\m5.addrM64 [35]), .A(n3432), .Z(n3003) );
  CANR1X1 U5909 ( .A(n3434), .B(\m0.addrM64 [35]), .C(n3003), .Z(n3004) );
  CND3X2 U5910 ( .A(n3006), .B(n3005), .C(n3004), .Z(n4173) );
  CAN2XL U5911 ( .A(\s6.addr [17]), .B(n4173), .Z(\s6.addr [35]) );
  CAN2XL U5912 ( .A(\s6.addr [17]), .B(n4165), .Z(\s6.addr [51]) );
  CAN2XL U5913 ( .A(\s6.addr [17]), .B(n4130), .Z(\s6.SbusIn [59]) );
  CIVX2 U5914 ( .A(\m5.addrM64 [43]), .Z(n3008) );
  CND2X1 U5915 ( .A(n3435), .B(\m6.addrM64 [43]), .Z(n3007) );
  COND1X1 U5916 ( .A(n3432), .B(n3008), .C(n3007), .Z(n3009) );
  CNR2X1 U5917 ( .A(n3010), .B(n3009), .Z(n3014) );
  CNR2IX1 U5918 ( .B(\m4.addrM64 [43]), .A(n3439), .Z(n3011) );
  CANR1X1 U5919 ( .A(n3431), .B(\m1.addrM64 [43]), .C(n3011), .Z(n3013) );
  CND2X2 U5920 ( .A(n3289), .B(\m3.addrM64 [43]), .Z(n3012) );
  CND3X2 U5921 ( .A(n3014), .B(n3013), .C(n3012), .Z(n4122) );
  CAN2XL U5922 ( .A(n4405), .B(n4122), .Z(\s5.addr [43]) );
  CAN2XL U5923 ( .A(n4405), .B(n4125), .Z(\s5.SbusIn [61]) );
  CIVX2 U5924 ( .A(n3473), .Z(n4231) );
  CNR2X1 U5925 ( .A(n2223), .B(n4231), .Z(\s8.SbusIn [22]) );
  CAN2XL U5926 ( .A(\s14.addr[18] ), .B(n4237), .Z(\s14.SbusIn [35]) );
  CND2XL U5927 ( .A(n3431), .B(\m1.DoutM [41]), .Z(n3016) );
  CND2XL U5928 ( .A(n3436), .B(\m2.DoutM [41]), .Z(n3015) );
  CND2X1 U5929 ( .A(n3016), .B(n3015), .Z(n3018) );
  CNR2IX1 U5930 ( .B(\m4.DoutM [41]), .A(n3439), .Z(n3017) );
  CNR2X1 U5931 ( .A(n3018), .B(n3017), .Z(n3022) );
  CANR2X1 U5932 ( .A(n3420), .B(\m3.DoutM [41]), .C(\m6.DoutM [41]), .D(n3435), 
        .Z(n3021) );
  CNR2IX1 U5933 ( .B(\m5.DoutM [41]), .A(n3432), .Z(n3019) );
  CANR1X1 U5934 ( .A(n3434), .B(\m0.DoutM [41]), .C(n3019), .Z(n3020) );
  CND3X2 U5935 ( .A(n3022), .B(n3021), .C(n3020), .Z(n4142) );
  CAN2XL U5936 ( .A(\s14.addr[18] ), .B(n4142), .Z(\s14.SbusIn [41]) );
  CAN2XL U5937 ( .A(\s14.addr[18] ), .B(n4180), .Z(\s14.SbusIn [18]) );
  CND2X1 U5938 ( .A(n3430), .B(\m3.DoutM [49]), .Z(n3025) );
  CND2X1 U5939 ( .A(n3434), .B(\m0.DoutM [49]), .Z(n3024) );
  CND2X1 U5940 ( .A(n3431), .B(\m1.DoutM [49]), .Z(n3023) );
  CAN3X2 U5941 ( .A(n3025), .B(n3024), .C(n3023), .Z(n3029) );
  CNR2X1 U5942 ( .A(n3027), .B(n3026), .Z(n3028) );
  CND2X2 U5943 ( .A(n3029), .B(n3028), .Z(n3480) );
  CAN2XL U5944 ( .A(\s14.addr[18] ), .B(n3480), .Z(\s14.SbusIn [49]) );
  CND2X1 U5945 ( .A(n3434), .B(\m0.DoutM [8]), .Z(n3031) );
  CND2XL U5946 ( .A(n3436), .B(\m2.DoutM [8]), .Z(n3030) );
  CND2X1 U5947 ( .A(n3031), .B(n3030), .Z(n3033) );
  CNR2X1 U5948 ( .A(n3033), .B(n3032), .Z(n3037) );
  CNR2IX1 U5949 ( .B(\m4.DoutM [8]), .A(n3439), .Z(n3034) );
  CANR1X1 U5950 ( .A(n3431), .B(\m1.DoutM [8]), .C(n3034), .Z(n3036) );
  CND2X1 U5951 ( .A(n3420), .B(\m3.DoutM [8]), .Z(n3035) );
  CND3X2 U5952 ( .A(n3037), .B(n3036), .C(n3035), .Z(n4116) );
  CAN2XL U5953 ( .A(\s14.addr[18] ), .B(n4116), .Z(\s14.SbusIn [8]) );
  CAN2XL U5954 ( .A(\s14.addr[18] ), .B(n4126), .Z(\s14.SbusIn [62]) );
  CIVX12 U5955 ( .A(n3453), .Z(\s1.addr [19]) );
  CIVX16 U5956 ( .A(n3378), .Z(\s10.addr [17]) );
  CIVX12 U5957 ( .A(n3038), .Z(\s11.addr[19] ) );
  CNR2XL U5958 ( .A(n3380), .B(n5587), .Z(\m0.MinData [63]) );
  CNR2XL U5959 ( .A(n3380), .B(n5570), .Z(\m0.MinData [47]) );
  CNR2XL U5960 ( .A(n3380), .B(n5585), .Z(\m0.MinData [61]) );
  CNR2XL U5961 ( .A(n3380), .B(n5571), .Z(\m0.MinData [48]) );
  CNR2XL U5962 ( .A(n3380), .B(n5568), .Z(\m0.MinData [45]) );
  CNR2XL U5963 ( .A(n3380), .B(n5584), .Z(\m0.MinData [60]) );
  CNR2XL U5964 ( .A(n3380), .B(n5569), .Z(\m0.MinData [46]) );
  CNR2XL U5965 ( .A(n3380), .B(n5586), .Z(\m0.MinData [62]) );
  CNR2XL U5966 ( .A(n3380), .B(n5572), .Z(\m0.MinData [49]) );
  CIVX3 U5967 ( .A(\m6.ack ), .Z(n3381) );
  CNR2XL U5968 ( .A(n3381), .B(n5568), .Z(\m6.MinData [45]) );
  CNR2XL U5969 ( .A(n3381), .B(n5569), .Z(\m6.MinData [46]) );
  CNR2XL U5970 ( .A(n3381), .B(n5570), .Z(\m6.MinData [47]) );
  CNR2XL U5971 ( .A(n3381), .B(n5571), .Z(\m6.MinData [48]) );
  CNR2XL U5972 ( .A(n3381), .B(n5572), .Z(\m6.MinData [49]) );
  CNR2XL U5973 ( .A(n3381), .B(n5584), .Z(\m6.MinData [60]) );
  CNR2XL U5974 ( .A(n3381), .B(n5585), .Z(\m6.MinData [61]) );
  CNR2XL U5975 ( .A(n3381), .B(n5586), .Z(\m6.MinData [62]) );
  CNR2XL U5976 ( .A(n3381), .B(n5587), .Z(\m6.MinData [63]) );
  CIVX2 U5977 ( .A(\m2.ack ), .Z(n3382) );
  CNR2XL U5978 ( .A(n3382), .B(n5574), .Z(\m2.MinData [50]) );
  CNR2XL U5979 ( .A(n3382), .B(n5575), .Z(\m2.MinData [51]) );
  CNR2XL U5980 ( .A(n3382), .B(n5576), .Z(\m2.MinData [52]) );
  CNR2XL U5981 ( .A(n3382), .B(n5577), .Z(\m2.MinData [53]) );
  CNR2XL U5982 ( .A(n3382), .B(n5578), .Z(\m2.MinData [54]) );
  CNR2XL U5983 ( .A(n3382), .B(n5584), .Z(\m2.MinData [60]) );
  CNR2XL U5984 ( .A(n3382), .B(n5585), .Z(\m2.MinData [61]) );
  CNR2XL U5985 ( .A(n3382), .B(n5586), .Z(\m2.MinData [62]) );
  CNR2XL U5986 ( .A(n3382), .B(n5587), .Z(\m2.MinData [63]) );
  CAN2X1 U5987 ( .A(\s4.en ), .B(n3478), .Z(\s4.addr [6]) );
  CAN2X1 U5988 ( .A(\s4.en ), .B(n4237), .Z(\s4.SbusIn [35]) );
  CIVX2 U5989 ( .A(n3459), .Z(n4333) );
  CAN2X1 U5990 ( .A(\s4.addr[14] ), .B(n4333), .Z(\s4.addr [3]) );
  CAN2X1 U5991 ( .A(\s4.en ), .B(n3456), .Z(\s4.addr [7]) );
  CAN2XL U5992 ( .A(\s8.addr[17] ), .B(n4141), .Z(\s8.SbusIn [25]) );
  CAN2XL U5993 ( .A(\s8.en ), .B(n3465), .Z(\s8.SbusIn [11]) );
  CAN2XL U5994 ( .A(\s8.addr[17] ), .B(n4192), .Z(\s8.SbusIn [2]) );
  CND2X1 U5995 ( .A(n3431), .B(\m1.DoutM [6]), .Z(n3040) );
  CND2XL U5996 ( .A(n3436), .B(\m2.DoutM [6]), .Z(n3039) );
  CND2X1 U5997 ( .A(n3040), .B(n3039), .Z(n3042) );
  CNR2IX1 U5998 ( .B(\m4.DoutM [6]), .A(n3439), .Z(n3041) );
  CNR2X1 U5999 ( .A(n3042), .B(n3041), .Z(n3046) );
  CANR2X1 U6000 ( .A(n3361), .B(\m3.DoutM [6]), .C(\m6.DoutM [6]), .D(n3435), 
        .Z(n3045) );
  CNR2IX1 U6001 ( .B(\m5.DoutM [6]), .A(n3432), .Z(n3043) );
  CANR1X1 U6002 ( .A(n3434), .B(\m0.DoutM [6]), .C(n3043), .Z(n3044) );
  CND3X2 U6003 ( .A(n3046), .B(n3045), .C(n3044), .Z(n4329) );
  CAN2XL U6004 ( .A(\s8.en ), .B(n4329), .Z(\s8.SbusIn [6]) );
  CIVX2 U6005 ( .A(n3477), .Z(n4244) );
  CNR2X1 U6006 ( .A(n3451), .B(n4244), .Z(\s7.addr [59]) );
  CIVDX3 U6007 ( .A(n3047), .Z0(n3468), .Z1(n4339) );
  CAN2X1 U6008 ( .A(\s7.addr[19] ), .B(n4339), .Z(\s7.addr [1]) );
  CND2XL U6009 ( .A(n3431), .B(\m1.addrM64 [57]), .Z(n3049) );
  CND2XL U6010 ( .A(n3436), .B(\m2.addrM64 [57]), .Z(n3048) );
  CND2X1 U6011 ( .A(n3049), .B(n3048), .Z(n3051) );
  CAN2XL U6012 ( .A(n3424), .B(\m4.addrM64 [57]), .Z(n3050) );
  CNR2X1 U6013 ( .A(n3051), .B(n3050), .Z(n3055) );
  CANR2X1 U6014 ( .A(n3420), .B(\m3.addrM64 [57]), .C(\m6.addrM64 [57]), .D(
        n3435), .Z(n3054) );
  CNR2IX1 U6015 ( .B(\m5.addrM64 [57]), .A(n3432), .Z(n3052) );
  CANR1X1 U6016 ( .A(n3434), .B(\m0.addrM64 [57]), .C(n3052), .Z(n3053) );
  CND3X2 U6017 ( .A(n3055), .B(n3054), .C(n3053), .Z(n4207) );
  CAN2XL U6018 ( .A(\s7.en ), .B(n4207), .Z(\s7.addr [57]) );
  CAN2XL U6019 ( .A(\s8.addr[17] ), .B(n4169), .Z(\s8.SbusIn [15]) );
  CND2X1 U6020 ( .A(n3371), .B(\m3.DoutM [5]), .Z(n3058) );
  CND2X1 U6021 ( .A(n3434), .B(\m0.DoutM [5]), .Z(n3057) );
  CND2X1 U6022 ( .A(n3431), .B(\m1.DoutM [5]), .Z(n3056) );
  CAN3X2 U6023 ( .A(n3058), .B(n3057), .C(n3056), .Z(n3066) );
  CIVX2 U6024 ( .A(\m5.DoutM [5]), .Z(n3060) );
  CND2X1 U6025 ( .A(n3435), .B(\m6.DoutM [5]), .Z(n3059) );
  CND2X1 U6026 ( .A(n3436), .B(\m2.DoutM [5]), .Z(n3062) );
  CND2XL U6027 ( .A(n3424), .B(\m4.DoutM [5]), .Z(n3061) );
  CND2X1 U6028 ( .A(n3062), .B(n3061), .Z(n3063) );
  CNR2X1 U6029 ( .A(n3064), .B(n3063), .Z(n3065) );
  CND2X2 U6030 ( .A(n3066), .B(n3065), .Z(n3469) );
  CAN2XL U6031 ( .A(\s12.addr[10] ), .B(n3469), .Z(\s12.SbusIn [5]) );
  CAN2XL U6032 ( .A(n4336), .B(n4242), .Z(\s7.addr [56]) );
  CAN2XL U6033 ( .A(\s8.addr[15] ), .B(n4121), .Z(\s8.SbusIn [48]) );
  CAN2XL U6034 ( .A(\s12.addr[10] ), .B(n4329), .Z(\s12.SbusIn [6]) );
  CAN2XL U6035 ( .A(\s8.en ), .B(n4171), .Z(\s8.SbusIn [32]) );
  CNIVX2 U6036 ( .A(n3451), .Z(n3452) );
  CND2XL U6037 ( .A(n3431), .B(\m1.addrM64 [41]), .Z(n3068) );
  CND2XL U6038 ( .A(n3436), .B(\m2.addrM64 [41]), .Z(n3067) );
  CND2X1 U6039 ( .A(n3068), .B(n3067), .Z(n3070) );
  CNR2IX1 U6040 ( .B(\m4.addrM64 [41]), .A(n3439), .Z(n3069) );
  CNR2X1 U6041 ( .A(n3070), .B(n3069), .Z(n3074) );
  CANR2X1 U6042 ( .A(n3137), .B(\m3.addrM64 [41]), .C(\m6.addrM64 [41]), .D(
        n3435), .Z(n3073) );
  CNR2IX1 U6043 ( .B(\m5.addrM64 [41]), .A(n3432), .Z(n3071) );
  CANR1X1 U6044 ( .A(n3434), .B(\m0.addrM64 [41]), .C(n3071), .Z(n3072) );
  CND3X2 U6045 ( .A(n3074), .B(n3073), .C(n3072), .Z(n3471) );
  CIVX2 U6046 ( .A(n3471), .Z(n4300) );
  CNR2X1 U6047 ( .A(n3452), .B(n4300), .Z(\s7.addr [41]) );
  CND2X1 U6048 ( .A(n3361), .B(\m3.DoutM [31]), .Z(n3077) );
  CND2X1 U6049 ( .A(n3434), .B(\m0.DoutM [31]), .Z(n3076) );
  CND2X1 U6050 ( .A(n3431), .B(\m1.DoutM [31]), .Z(n3075) );
  CAN3X2 U6051 ( .A(n3077), .B(n3076), .C(n3075), .Z(n3083) );
  CIVX2 U6052 ( .A(\m5.DoutM [31]), .Z(n3079) );
  CND2X1 U6053 ( .A(n3435), .B(\m6.DoutM [31]), .Z(n3078) );
  CNR2X1 U6054 ( .A(n3081), .B(n3080), .Z(n3082) );
  CND2X2 U6055 ( .A(n3083), .B(n3082), .Z(n4119) );
  CAN2XL U6056 ( .A(\s8.en ), .B(n4119), .Z(\s8.SbusIn [31]) );
  CND2X1 U6057 ( .A(n3434), .B(\m0.addrM64 [39]), .Z(n3085) );
  CND2XL U6058 ( .A(n3436), .B(\m2.addrM64 [39]), .Z(n3084) );
  CND2X1 U6059 ( .A(n3085), .B(n3084), .Z(n3089) );
  CIVX2 U6060 ( .A(\m5.addrM64 [39]), .Z(n3087) );
  CND2X1 U6061 ( .A(n3435), .B(\m6.addrM64 [39]), .Z(n3086) );
  CNR2X1 U6062 ( .A(n3089), .B(n3088), .Z(n3094) );
  CANR2X1 U6063 ( .A(n3431), .B(\m1.addrM64 [39]), .C(\m3.addrM64 [39]), .D(
        n3090), .Z(n3093) );
  CNR2IX1 U6064 ( .B(\m4.addrM64 [39]), .A(n3439), .Z(n3091) );
  CIVX2 U6065 ( .A(n3091), .Z(n3092) );
  CAN2XL U6066 ( .A(\s7.en ), .B(n4177), .Z(\s7.addr [39]) );
  CND2X1 U6067 ( .A(n3434), .B(\m0.addrM64 [38]), .Z(n3096) );
  CND2XL U6068 ( .A(n3436), .B(\m2.addrM64 [38]), .Z(n3095) );
  CND2X1 U6069 ( .A(n3096), .B(n3095), .Z(n3098) );
  CNR2X1 U6070 ( .A(n3098), .B(n3097), .Z(n3102) );
  CNR2IX1 U6071 ( .B(\m4.addrM64 [38]), .A(n3439), .Z(n3099) );
  CANR1X1 U6072 ( .A(n3431), .B(\m1.addrM64 [38]), .C(n3099), .Z(n3101) );
  CND2X1 U6073 ( .A(n3361), .B(\m3.addrM64 [38]), .Z(n3100) );
  CND3X2 U6074 ( .A(n3102), .B(n3101), .C(n3100), .Z(n4204) );
  CAN2XL U6075 ( .A(\s7.addr[16] ), .B(n4204), .Z(\s7.addr [38]) );
  CAN2XL U6076 ( .A(\s8.addr[15] ), .B(n4178), .Z(\s8.SbusIn [34]) );
  CND2XL U6077 ( .A(n3431), .B(\m1.addrM64 [37]), .Z(n3104) );
  CND2XL U6078 ( .A(n3436), .B(\m2.addrM64 [37]), .Z(n3103) );
  CND2X1 U6079 ( .A(n3104), .B(n3103), .Z(n3106) );
  CNR2IX1 U6080 ( .B(\m4.addrM64 [37]), .A(n3439), .Z(n3105) );
  CNR2X1 U6081 ( .A(n3106), .B(n3105), .Z(n3110) );
  CANR2X1 U6082 ( .A(n3420), .B(\m3.addrM64 [37]), .C(\m6.addrM64 [37]), .D(
        n3435), .Z(n3109) );
  CNR2IX1 U6083 ( .B(\m5.addrM64 [37]), .A(n3432), .Z(n3107) );
  CANR1X1 U6084 ( .A(n3434), .B(\m0.addrM64 [37]), .C(n3107), .Z(n3108) );
  CND3X2 U6085 ( .A(n3110), .B(n3109), .C(n3108), .Z(n3464) );
  CAN2XL U6086 ( .A(\s7.addr[19] ), .B(n3464), .Z(\s7.addr [37]) );
  CAN2XL U6087 ( .A(\s8.en ), .B(n4158), .Z(\s8.SbusIn [21]) );
  CAN2X1 U6088 ( .A(\s8.addr[17] ), .B(n4237), .Z(\s8.SbusIn [35]) );
  CAN2XL U6089 ( .A(\s7.addr[19] ), .B(n4160), .Z(\s7.addr [31]) );
  CAN2XL U6090 ( .A(\s8.en ), .B(n4116), .Z(\s8.SbusIn [8]) );
  CAN2XL U6091 ( .A(\s8.addr[17] ), .B(n4185), .Z(\s8.SbusIn [0]) );
  CAN2XL U6092 ( .A(\s8.en ), .B(n4190), .Z(\s8.SbusIn [1]) );
  CND2XL U6093 ( .A(n3434), .B(\m0.DoutM [37]), .Z(n3112) );
  CND2X1 U6094 ( .A(n3436), .B(\m2.DoutM [37]), .Z(n3111) );
  CND2X1 U6095 ( .A(n3112), .B(n3111), .Z(n3116) );
  CIVX2 U6096 ( .A(\m5.DoutM [37]), .Z(n3114) );
  CND2X1 U6097 ( .A(n3435), .B(\m6.DoutM [37]), .Z(n3113) );
  COND1X1 U6098 ( .A(n3432), .B(n3114), .C(n3113), .Z(n3115) );
  CNR2X1 U6099 ( .A(n3116), .B(n3115), .Z(n3120) );
  CANR2X1 U6100 ( .A(n3431), .B(\m1.DoutM [37]), .C(\m3.DoutM [37]), .D(n3137), 
        .Z(n3119) );
  CNR2IX1 U6101 ( .B(\m4.DoutM [37]), .A(n3439), .Z(n3117) );
  CIVX2 U6102 ( .A(n3117), .Z(n3118) );
  CND3X2 U6103 ( .A(n3120), .B(n3119), .C(n3118), .Z(n4196) );
  CAN2XL U6104 ( .A(\s8.addr[15] ), .B(n4196), .Z(\s8.SbusIn [37]) );
  CIVX2 U6105 ( .A(n3467), .Z(n4246) );
  CNR2X1 U6106 ( .A(n3452), .B(n4246), .Z(\s7.addr [27]) );
  CAN2XL U6107 ( .A(\s8.addr[15] ), .B(n4193), .Z(\s8.SbusIn [9]) );
  CAN2XL U6108 ( .A(\s8.addr[15] ), .B(n4197), .Z(\s8.SbusIn [29]) );
  CND2X1 U6109 ( .A(n3434), .B(\m0.addrM64 [50]), .Z(n3122) );
  CND2XL U6110 ( .A(n3436), .B(\m2.addrM64 [50]), .Z(n3121) );
  CND2X1 U6111 ( .A(n3122), .B(n3121), .Z(n3126) );
  CIVX2 U6112 ( .A(\m5.addrM64 [50]), .Z(n3124) );
  CND2X1 U6113 ( .A(n3435), .B(\m6.addrM64 [50]), .Z(n3123) );
  CNR2X1 U6114 ( .A(n3126), .B(n3125), .Z(n3130) );
  CANR2X1 U6115 ( .A(n3431), .B(\m1.addrM64 [50]), .C(\m3.addrM64 [50]), .D(
        n3420), .Z(n3129) );
  CNR2IX1 U6116 ( .B(\m4.addrM64 [50]), .A(n3439), .Z(n3127) );
  CIVX2 U6117 ( .A(n3127), .Z(n3128) );
  CAN2XL U6118 ( .A(\s7.en ), .B(n4164), .Z(\s7.addr [50]) );
  CND2X1 U6119 ( .A(n3434), .B(\m0.addrM64 [23]), .Z(n3132) );
  CND2X1 U6120 ( .A(n3436), .B(\m2.addrM64 [23]), .Z(n3131) );
  CND2X1 U6121 ( .A(n3132), .B(n3131), .Z(n3136) );
  CIVX2 U6122 ( .A(\m5.addrM64 [23]), .Z(n3134) );
  CND2X1 U6123 ( .A(n3435), .B(\m6.addrM64 [23]), .Z(n3133) );
  CNR2X1 U6124 ( .A(n3136), .B(n3135), .Z(n3141) );
  CANR2X1 U6125 ( .A(n3431), .B(\m1.addrM64 [23]), .C(\m3.addrM64 [23]), .D(
        n3137), .Z(n3140) );
  CNR2IX1 U6126 ( .B(\m4.addrM64 [23]), .A(n3439), .Z(n3138) );
  CIVX2 U6127 ( .A(n3138), .Z(n3139) );
  CAN2XL U6128 ( .A(n4336), .B(n4118), .Z(\s7.addr [23]) );
  CND2XL U6129 ( .A(n3431), .B(\m1.addrM64 [60]), .Z(n3143) );
  CND2XL U6130 ( .A(n3436), .B(\m2.addrM64 [60]), .Z(n3142) );
  CND2X1 U6131 ( .A(n3143), .B(n3142), .Z(n3145) );
  CAN2XL U6132 ( .A(n3424), .B(\m4.addrM64 [60]), .Z(n3144) );
  CNR2X1 U6133 ( .A(n3145), .B(n3144), .Z(n3149) );
  CANR2X1 U6134 ( .A(n3361), .B(\m3.addrM64 [60]), .C(\m6.addrM64 [60]), .D(
        n3435), .Z(n3148) );
  CNR2IX1 U6135 ( .B(\m5.addrM64 [60]), .A(n3432), .Z(n3146) );
  CANR1X1 U6136 ( .A(n3434), .B(\m0.addrM64 [60]), .C(n3146), .Z(n3147) );
  CND3X2 U6137 ( .A(n3149), .B(n3148), .C(n3147), .Z(n3482) );
  CAN2XL U6138 ( .A(\s7.addr[16] ), .B(n3482), .Z(\s7.addr [60]) );
  CNR2X1 U6139 ( .A(n3151), .B(n3150), .Z(n3155) );
  CANR2X1 U6140 ( .A(n3431), .B(\m1.DoutM [14]), .C(\m3.DoutM [14]), .D(n3420), 
        .Z(n3154) );
  CNR2IX1 U6141 ( .B(\m4.DoutM [14]), .A(n3439), .Z(n3152) );
  CIVX2 U6142 ( .A(n3152), .Z(n3153) );
  CND3X2 U6143 ( .A(n3155), .B(n3154), .C(n3153), .Z(n3474) );
  CAN2X1 U6144 ( .A(\s8.addr[17] ), .B(n3474), .Z(\s8.SbusIn [14]) );
  CAN2X1 U6145 ( .A(\s8.en ), .B(n4173), .Z(\s8.addr [35]) );
  CND2XL U6146 ( .A(n3431), .B(\m1.addrM64 [58]), .Z(n3157) );
  CND2XL U6147 ( .A(n3436), .B(\m2.addrM64 [58]), .Z(n3156) );
  CND2X1 U6148 ( .A(n3157), .B(n3156), .Z(n3159) );
  CAN2XL U6149 ( .A(n3424), .B(\m4.addrM64 [58]), .Z(n3158) );
  CNR2X1 U6150 ( .A(n3159), .B(n3158), .Z(n3163) );
  CANR2X1 U6151 ( .A(n3420), .B(\m3.addrM64 [58]), .C(\m6.addrM64 [58]), .D(
        n3435), .Z(n3162) );
  CNR2IX1 U6152 ( .B(\m5.addrM64 [58]), .A(n3432), .Z(n3160) );
  CANR1X1 U6153 ( .A(n3434), .B(\m0.addrM64 [58]), .C(n3160), .Z(n3161) );
  CND3X2 U6154 ( .A(n3163), .B(n3162), .C(n3161), .Z(n4202) );
  CAN2XL U6155 ( .A(\s8.addr[15] ), .B(n4202), .Z(\s8.addr [58]) );
  CAN2XL U6156 ( .A(\s8.en ), .B(n4179), .Z(\s8.addr [33]) );
  CAN2XL U6157 ( .A(\s8.addr[15] ), .B(n4151), .Z(\s8.addr [61]) );
  CAN2XL U6158 ( .A(\s8.addr[15] ), .B(n3479), .Z(\s8.addr [62]) );
  CND2X1 U6159 ( .A(n3431), .B(\m1.DoutM [42]), .Z(n3165) );
  CND2XL U6160 ( .A(n3436), .B(\m2.DoutM [42]), .Z(n3164) );
  CND2X1 U6161 ( .A(n3165), .B(n3164), .Z(n3167) );
  CNR2IX1 U6162 ( .B(\m4.DoutM [42]), .A(n3439), .Z(n3166) );
  CNR2X1 U6163 ( .A(n3167), .B(n3166), .Z(n3171) );
  CANR2X1 U6164 ( .A(n3420), .B(\m3.DoutM [42]), .C(\m6.DoutM [42]), .D(n3435), 
        .Z(n3170) );
  CNR2IX1 U6165 ( .B(\m5.DoutM [42]), .A(n3432), .Z(n3168) );
  CANR1X1 U6166 ( .A(n3434), .B(\m0.DoutM [42]), .C(n3168), .Z(n3169) );
  CND3X2 U6167 ( .A(n3171), .B(n3170), .C(n3169), .Z(n4144) );
  CAN2XL U6168 ( .A(\s12.addr[10] ), .B(n4144), .Z(\s12.SbusIn [42]) );
  CAN2XL U6169 ( .A(\s8.en ), .B(n3467), .Z(\s8.addr [27]) );
  CAN2X1 U6170 ( .A(\s12.addr[10] ), .B(n4333), .Z(\s12.addr [3]) );
  CAN2XL U6171 ( .A(\s8.en ), .B(n4136), .Z(\s8.addr [46]) );
  CAN2X1 U6172 ( .A(\s12.addr[10] ), .B(n4339), .Z(\s12.addr [1]) );
  CAN2XL U6173 ( .A(\s8.en ), .B(n4137), .Z(\s8.addr [48]) );
  CAN2XL U6174 ( .A(\s8.en ), .B(n4164), .Z(\s8.addr [50]) );
  CAN2XL U6175 ( .A(\s8.addr[15] ), .B(n4122), .Z(\s8.addr [43]) );
  CANR2X1 U6176 ( .A(n3431), .B(\m1.addrM64 [42]), .C(\m3.addrM64 [42]), .D(
        n3299), .Z(n3179) );
  CNR2IX1 U6177 ( .B(\m5.addrM64 [42]), .A(n3432), .Z(n3172) );
  CND2XL U6178 ( .A(n3435), .B(\m6.addrM64 [42]), .Z(n3174) );
  CND2X1 U6179 ( .A(n3436), .B(\m2.addrM64 [42]), .Z(n3173) );
  CND2X1 U6180 ( .A(n3174), .B(n3173), .Z(n3176) );
  CNR2IX1 U6181 ( .B(\m4.addrM64 [42]), .A(n3439), .Z(n3175) );
  CNR2X1 U6182 ( .A(n3176), .B(n3175), .Z(n3177) );
  CND3X2 U6183 ( .A(n3179), .B(n3178), .C(n3177), .Z(n4153) );
  CAN2XL U6184 ( .A(\s8.en ), .B(n4153), .Z(\s8.addr [42]) );
  CAN2X1 U6185 ( .A(n3420), .B(\m3.addrM64 [52]), .Z(n3180) );
  CND2X1 U6186 ( .A(n3434), .B(\m0.addrM64 [52]), .Z(n3182) );
  CNR2IX1 U6187 ( .B(\m5.addrM64 [52]), .A(n3432), .Z(n3181) );
  CNR2IX1 U6188 ( .B(n3182), .A(n3181), .Z(n3186) );
  CAN2XL U6189 ( .A(n3424), .B(\m4.addrM64 [52]), .Z(n3183) );
  CNR2X1 U6190 ( .A(n3184), .B(n3183), .Z(n3185) );
  CND3X2 U6191 ( .A(n3187), .B(n3186), .C(n3185), .Z(n4166) );
  CAN2X1 U6192 ( .A(\s8.en ), .B(n4166), .Z(\s8.addr [52]) );
  CANR2X1 U6193 ( .A(n3431), .B(\m1.DoutM [54]), .C(\m3.DoutM [54]), .D(n3420), 
        .Z(n3195) );
  CNR2IX1 U6194 ( .B(\m5.DoutM [54]), .A(n3432), .Z(n3188) );
  CANR1X1 U6195 ( .A(n3434), .B(\m0.DoutM [54]), .C(n3188), .Z(n3194) );
  CND2XL U6196 ( .A(n3435), .B(\m6.DoutM [54]), .Z(n3190) );
  CND2X1 U6197 ( .A(n3436), .B(\m2.DoutM [54]), .Z(n3189) );
  CND2X1 U6198 ( .A(n3190), .B(n3189), .Z(n3192) );
  CNR2IX1 U6199 ( .B(\m4.DoutM [54]), .A(n3439), .Z(n3191) );
  CNR2X1 U6200 ( .A(n3192), .B(n3191), .Z(n3193) );
  CND3X2 U6201 ( .A(n3195), .B(n3194), .C(n3193), .Z(n4175) );
  CAN2XL U6202 ( .A(\s12.addr[10] ), .B(n4175), .Z(\s12.SbusIn [54]) );
  CAN2XL U6203 ( .A(\s8.en ), .B(n4177), .Z(\s8.addr [39]) );
  CAN2XL U6204 ( .A(\s8.en ), .B(n4148), .Z(\s8.addr [54]) );
  CAN2XL U6205 ( .A(\s12.addr[10] ), .B(n4163), .Z(\s12.SbusIn [51]) );
  CAN2XL U6206 ( .A(\s8.addr[17] ), .B(n4124), .Z(\s8.addr [36]) );
  CAN2XL U6207 ( .A(\s8.en ), .B(n4126), .Z(\s8.SbusIn [62]) );
  CAN2XL U6208 ( .A(\s7.addr[16] ), .B(n4178), .Z(\s7.SbusIn [34]) );
  CAN2XL U6209 ( .A(\s8.en ), .B(n4167), .Z(\s8.SbusIn [60]) );
  CAN2XL U6210 ( .A(n4336), .B(n4215), .Z(\s7.SbusIn [36]) );
  CAN2X1 U6211 ( .A(n3420), .B(\m3.DoutM [58]), .Z(n3196) );
  CNR2IX1 U6212 ( .B(\m5.DoutM [58]), .A(n3432), .Z(n3197) );
  CNR2IX1 U6213 ( .B(\m4.DoutM [58]), .A(n3439), .Z(n3198) );
  CNR2X1 U6214 ( .A(n3199), .B(n3198), .Z(n3200) );
  CND3X2 U6215 ( .A(n3202), .B(n3201), .C(n3200), .Z(n4168) );
  CAN2XL U6216 ( .A(\s8.addr[15] ), .B(n4168), .Z(\s8.SbusIn [58]) );
  CAN2XL U6217 ( .A(\s7.en ), .B(n4142), .Z(\s7.SbusIn [41]) );
  CAN2XL U6218 ( .A(\s12.addr[10] ), .B(n3465), .Z(\s12.SbusIn [11]) );
  CAN2XL U6219 ( .A(\s8.en ), .B(n4175), .Z(\s8.SbusIn [54]) );
  CAN2XL U6220 ( .A(\s8.en ), .B(n4170), .Z(\s8.SbusIn [53]) );
  CAN2XL U6221 ( .A(\s8.addr[15] ), .B(n4163), .Z(\s8.SbusIn [51]) );
  CAN2XL U6222 ( .A(\s8.en ), .B(n4127), .Z(\s8.SbusIn [50]) );
  CND2X1 U6223 ( .A(n3434), .B(\m0.DoutM [55]), .Z(n3204) );
  CND2XL U6224 ( .A(n3436), .B(\m2.DoutM [55]), .Z(n3203) );
  CIVX2 U6225 ( .A(\m5.DoutM [55]), .Z(n3206) );
  CND2X1 U6226 ( .A(n3435), .B(\m6.DoutM [55]), .Z(n3205) );
  CAN2XL U6227 ( .A(\s7.en ), .B(n3461), .Z(\s7.SbusIn [55]) );
  CAN2X1 U6228 ( .A(\s12.addr[10] ), .B(n4201), .Z(\s12.addr [55]) );
  CAN2XL U6229 ( .A(\s7.addr[19] ), .B(n4200), .Z(\s7.SbusIn [3]) );
  CAN2XL U6230 ( .A(\s7.addr[16] ), .B(n4193), .Z(\s7.SbusIn [9]) );
  CAN2XL U6231 ( .A(n4336), .B(n3481), .Z(\s7.SbusIn [12]) );
  CIVX1 U6232 ( .A(n3454), .Z(n3455) );
  CAN2X1 U6233 ( .A(\s8.addr[17] ), .B(n3455), .Z(\s8.addr [9]) );
  CND2XL U6234 ( .A(n3431), .B(\m1.DoutM [17]), .Z(n3208) );
  CND2XL U6235 ( .A(n3436), .B(\m2.DoutM [17]), .Z(n3207) );
  CND2X1 U6236 ( .A(n3208), .B(n3207), .Z(n3210) );
  CNR2IX1 U6237 ( .B(\m4.DoutM [17]), .A(n3439), .Z(n3209) );
  CNR2X1 U6238 ( .A(n3210), .B(n3209), .Z(n3214) );
  CANR2X1 U6239 ( .A(n3299), .B(\m3.DoutM [17]), .C(\m6.DoutM [17]), .D(n3435), 
        .Z(n3213) );
  CNR2IX1 U6240 ( .B(\m5.DoutM [17]), .A(n3432), .Z(n3211) );
  CANR1X1 U6241 ( .A(n3434), .B(\m0.DoutM [17]), .C(n3211), .Z(n3212) );
  CND3X2 U6242 ( .A(n3214), .B(n3213), .C(n3212), .Z(n4172) );
  CAN2XL U6243 ( .A(\s7.en ), .B(n4172), .Z(\s7.SbusIn [17]) );
  CAN2X1 U6244 ( .A(\s8.addr[17] ), .B(n4333), .Z(\s8.addr [3]) );
  CAN2XL U6245 ( .A(n5445), .B(n3469), .Z(\s5.SbusIn [5]) );
  CAN2XL U6246 ( .A(n1844), .B(n4154), .Z(\s5.SbusIn [7]) );
  CANR2X1 U6247 ( .A(n3431), .B(\m1.DoutM [63]), .C(\m3.DoutM [63]), .D(n3420), 
        .Z(n3222) );
  CNR2IX1 U6248 ( .B(\m5.DoutM [63]), .A(n3432), .Z(n3215) );
  CND2X1 U6249 ( .A(n3435), .B(\m6.DoutM [63]), .Z(n3217) );
  CND2X1 U6250 ( .A(n3436), .B(\m2.DoutM [63]), .Z(n3216) );
  CND2X1 U6251 ( .A(n3217), .B(n3216), .Z(n3219) );
  CNR2IX1 U6252 ( .B(\m4.DoutM [63]), .A(n3439), .Z(n3218) );
  CNR2X1 U6253 ( .A(n3219), .B(n3218), .Z(n3220) );
  CND3X2 U6254 ( .A(n3222), .B(n3221), .C(n3220), .Z(n4120) );
  CAN2XL U6255 ( .A(n5445), .B(n4120), .Z(\s5.SbusIn [63]) );
  CAN2XL U6256 ( .A(n1844), .B(n4193), .Z(\s5.SbusIn [9]) );
  CAN2XL U6257 ( .A(n5445), .B(n4115), .Z(\s5.SbusIn [10]) );
  CAN2XL U6258 ( .A(n1844), .B(n3474), .Z(\s5.SbusIn [14]) );
  CAN2XL U6259 ( .A(n5445), .B(n4169), .Z(\s5.SbusIn [15]) );
  CAN2X1 U6260 ( .A(n3413), .B(n4405), .Z(\s5.addr [7]) );
  CAN2XL U6261 ( .A(n4405), .B(n4185), .Z(\s5.SbusIn [0]) );
  CAN2XL U6262 ( .A(n4405), .B(n4192), .Z(\s5.SbusIn [2]) );
  CAN2XL U6263 ( .A(n4405), .B(n4200), .Z(\s5.SbusIn [3]) );
  CAN2XL U6264 ( .A(n1844), .B(n4243), .Z(\s5.SbusIn [4]) );
  CAN2XL U6265 ( .A(n4405), .B(n4121), .Z(\s5.SbusIn [48]) );
  CAN2XL U6266 ( .A(n5445), .B(n4141), .Z(\s5.SbusIn [25]) );
  CAN2XL U6267 ( .A(n4405), .B(n4147), .Z(\s5.SbusIn [26]) );
  CAN2XL U6268 ( .A(n1844), .B(n3464), .Z(\s5.addr [37]) );
  CAN2XL U6269 ( .A(n5445), .B(n4117), .Z(\s5.SbusIn [28]) );
  CAN2XL U6270 ( .A(n4405), .B(n4145), .Z(\s5.SbusIn [30]) );
  CAN2XL U6271 ( .A(n4405), .B(n4119), .Z(\s5.SbusIn [31]) );
  CAN2XL U6272 ( .A(n4405), .B(n4171), .Z(\s5.SbusIn [32]) );
  CND2X1 U6273 ( .A(n3431), .B(\m1.DoutM [43]), .Z(n3224) );
  CND2XL U6274 ( .A(n3436), .B(\m2.DoutM [43]), .Z(n3223) );
  CND2X1 U6275 ( .A(n3224), .B(n3223), .Z(n3226) );
  CNR2IX1 U6276 ( .B(\m4.DoutM [43]), .A(n3439), .Z(n3225) );
  CNR2X1 U6277 ( .A(n3226), .B(n3225), .Z(n3230) );
  CANR2X1 U6278 ( .A(n3430), .B(\m3.DoutM [43]), .C(\m6.DoutM [43]), .D(n3435), 
        .Z(n3229) );
  CNR2IX1 U6279 ( .B(\m5.DoutM [43]), .A(n3432), .Z(n3227) );
  CND3X2 U6280 ( .A(n3230), .B(n3229), .C(n3228), .Z(n4132) );
  CAN2XL U6281 ( .A(n4405), .B(n4132), .Z(\s5.SbusIn [43]) );
  CAN2XL U6282 ( .A(n4405), .B(n4144), .Z(\s5.SbusIn [42]) );
  CAN2XL U6283 ( .A(n4405), .B(n4215), .Z(\s5.SbusIn [36]) );
  CIVX2 U6284 ( .A(\m5.DoutM [38]), .Z(n3233) );
  CND2XL U6285 ( .A(n3231), .B(\m6.DoutM [38]), .Z(n3232) );
  CNR2X1 U6286 ( .A(n3235), .B(n3234), .Z(n3239) );
  CANR2X1 U6287 ( .A(n3431), .B(\m1.DoutM [38]), .C(\m3.DoutM [38]), .D(n3361), 
        .Z(n3238) );
  CNR2IX1 U6288 ( .B(\m4.DoutM [38]), .A(n3439), .Z(n3236) );
  CIVX2 U6289 ( .A(n3236), .Z(n3237) );
  CND3X2 U6290 ( .A(n3239), .B(n3238), .C(n3237), .Z(n4232) );
  CAN2XL U6291 ( .A(n1844), .B(n4232), .Z(\s5.SbusIn [38]) );
  CAN2XL U6292 ( .A(n5445), .B(n4135), .Z(\s5.SbusIn [39]) );
  CAN2XL U6293 ( .A(n4405), .B(n4175), .Z(\s5.SbusIn [54]) );
  CAN2XL U6294 ( .A(n4405), .B(n3471), .Z(\s5.addr [41]) );
  CND2X1 U6295 ( .A(n3434), .B(\m0.addrM64 [24]), .Z(n3242) );
  CND2XL U6296 ( .A(n3436), .B(\m2.addrM64 [24]), .Z(n3241) );
  CND2X1 U6297 ( .A(n3242), .B(n3241), .Z(n3246) );
  CIVX2 U6298 ( .A(\m5.addrM64 [24]), .Z(n3244) );
  CND2X1 U6299 ( .A(n3435), .B(\m6.addrM64 [24]), .Z(n3243) );
  CNR2X1 U6300 ( .A(n3246), .B(n3245), .Z(n3250) );
  CANR2X1 U6301 ( .A(n3431), .B(\m1.addrM64 [24]), .C(\m3.addrM64 [24]), .D(
        n3420), .Z(n3249) );
  CNR2IX1 U6302 ( .B(\m4.addrM64 [24]), .A(n3439), .Z(n3247) );
  CIVX2 U6303 ( .A(n3247), .Z(n3248) );
  CAN2XL U6304 ( .A(n4405), .B(n4199), .Z(\s5.addr [24]) );
  CAN2XL U6305 ( .A(n4405), .B(n4158), .Z(\s5.SbusIn [21]) );
  CAN2XL U6306 ( .A(n1844), .B(n4204), .Z(\s5.addr [38]) );
  CAN2XL U6307 ( .A(n5445), .B(n4127), .Z(\s5.SbusIn [50]) );
  CAN2XL U6308 ( .A(\s6.addr [17]), .B(n4172), .Z(\s6.SbusIn [17]) );
  CAN2X1 U6309 ( .A(\s3.addr[14] ), .B(n4237), .Z(\s3.SbusIn [35]) );
  CAN2XL U6310 ( .A(\s6.addr [17]), .B(n4115), .Z(\s6.SbusIn [10]) );
  CND2XL U6311 ( .A(n3431), .B(\m1.DoutM [40]), .Z(n3253) );
  CND2XL U6312 ( .A(n3436), .B(\m2.DoutM [40]), .Z(n3252) );
  CND2X1 U6313 ( .A(n3253), .B(n3252), .Z(n3255) );
  CNR2IX1 U6314 ( .B(\m4.DoutM [40]), .A(n3439), .Z(n3254) );
  CNR2X1 U6315 ( .A(n3255), .B(n3254), .Z(n3259) );
  CANR2X1 U6316 ( .A(n3289), .B(\m3.DoutM [40]), .C(\m6.DoutM [40]), .D(n3435), 
        .Z(n3258) );
  CNR2IX1 U6317 ( .B(\m5.DoutM [40]), .A(n3432), .Z(n3256) );
  CANR1X1 U6318 ( .A(n3434), .B(\m0.DoutM [40]), .C(n3256), .Z(n3257) );
  CND3X2 U6319 ( .A(n3259), .B(n3258), .C(n3257), .Z(n4143) );
  CAN2XL U6320 ( .A(\s3.addr[14] ), .B(n4143), .Z(\s3.SbusIn [40]) );
  CAN2XL U6321 ( .A(\s6.addr [17]), .B(n4119), .Z(\s6.SbusIn [31]) );
  CAN2XL U6322 ( .A(\s6.addr [17]), .B(n3474), .Z(\s6.SbusIn [14]) );
  CNR2IX1 U6323 ( .B(\m5.DoutM [16]), .A(n3432), .Z(n3260) );
  CNR2IX1 U6324 ( .B(\m4.DoutM [16]), .A(n3439), .Z(n3261) );
  CIVX2 U6325 ( .A(n3261), .Z(n3264) );
  CANR2X1 U6326 ( .A(n3289), .B(\m3.DoutM [16]), .C(\m6.DoutM [16]), .D(n3435), 
        .Z(n3263) );
  CANR2X1 U6327 ( .A(n3434), .B(\m0.DoutM [16]), .C(n3436), .D(\m2.DoutM [16]), 
        .Z(n3262) );
  CND4X2 U6328 ( .A(n3265), .B(n3264), .C(n3263), .D(n3262), .Z(n3487) );
  CAN2XL U6329 ( .A(\s6.addr [17]), .B(n3487), .Z(\s6.SbusIn [16]) );
  CAN2XL U6330 ( .A(\s6.addr [17]), .B(n4152), .Z(\s6.SbusIn [19]) );
  CND2X1 U6331 ( .A(n3434), .B(\m0.addrM64 [53]), .Z(n3267) );
  CND2XL U6332 ( .A(n3436), .B(\m2.addrM64 [53]), .Z(n3266) );
  CND2X1 U6333 ( .A(n3267), .B(n3266), .Z(n3271) );
  CIVX2 U6334 ( .A(\m5.addrM64 [53]), .Z(n3269) );
  CND2X1 U6335 ( .A(n3435), .B(\m6.addrM64 [53]), .Z(n3268) );
  CNR2X1 U6336 ( .A(n3271), .B(n3270), .Z(n3275) );
  CAN2X1 U6337 ( .A(n3424), .B(\m4.addrM64 [53]), .Z(n3272) );
  CAN2XL U6338 ( .A(\s6.addr [17]), .B(n4174), .Z(\s6.addr [53]) );
  CAN2X1 U6339 ( .A(\s9.addr[16] ), .B(n4339), .Z(\s9.addr [1]) );
  CIVX8 U6340 ( .A(n3298), .Z(\s9.en ) );
  CAN2X1 U6341 ( .A(\s9.addr[7] ), .B(n4333), .Z(\s9.addr [3]) );
  CNR2IX1 U6342 ( .B(\m5.addrM64 [22]), .A(n3432), .Z(n3276) );
  CNR2IX1 U6343 ( .B(\m4.addrM64 [22]), .A(n3439), .Z(n3277) );
  CIVX2 U6344 ( .A(n3277), .Z(n3280) );
  CANR2X1 U6345 ( .A(n3435), .B(\m6.addrM64 [22]), .C(\m3.addrM64 [22]), .D(
        n3371), .Z(n3279) );
  CANR2X1 U6346 ( .A(n3434), .B(\m0.addrM64 [22]), .C(n3436), .D(
        \m2.addrM64 [22]), .Z(n3278) );
  CND4X2 U6347 ( .A(n3281), .B(n3280), .C(n3279), .D(n3278), .Z(n3462) );
  CAN2XL U6348 ( .A(\s9.addr[8] ), .B(n3462), .Z(\s9.addr [22]) );
  CAN2XL U6349 ( .A(\s3.addr[14] ), .B(n4200), .Z(\s3.SbusIn [3]) );
  CANR2X1 U6350 ( .A(n3431), .B(\m1.addrM64 [32]), .C(\m3.addrM64 [32]), .D(
        n3420), .Z(n3288) );
  CND2X1 U6351 ( .A(n3434), .B(\m0.addrM64 [32]), .Z(n3283) );
  CNR2IX1 U6352 ( .B(\m5.addrM64 [32]), .A(n3432), .Z(n3282) );
  CNR2IX1 U6353 ( .B(n3283), .A(n3282), .Z(n3287) );
  CNR2IX1 U6354 ( .B(\m4.addrM64 [32]), .A(n3439), .Z(n3284) );
  CNR2X1 U6355 ( .A(n3285), .B(n3284), .Z(n3286) );
  CND3X2 U6356 ( .A(n3288), .B(n3287), .C(n3286), .Z(n4157) );
  CAN2XL U6357 ( .A(\s3.addr[14] ), .B(n4157), .Z(\s3.addr [32]) );
  CAN2XL U6358 ( .A(\s9.addr[16] ), .B(n3467), .Z(\s9.addr [27]) );
  CAN2XL U6359 ( .A(\s9.addr[8] ), .B(n3479), .Z(\s9.addr [62]) );
  CIVX2 U6360 ( .A(n3482), .Z(n4251) );
  CNR2X1 U6361 ( .A(n3298), .B(n4251), .Z(\s9.addr [60]) );
  CNR2X1 U6362 ( .A(n3298), .B(n4244), .Z(\s9.addr [59]) );
  CAN2XL U6363 ( .A(\s9.addr[7] ), .B(n4207), .Z(\s9.addr [57]) );
  CAN2XL U6364 ( .A(\s9.addr[16] ), .B(n4242), .Z(\s9.addr [56]) );
  CIVX8 U6365 ( .A(n3298), .Z(n5590) );
  CAN2XL U6366 ( .A(\s9.addr[8] ), .B(n4201), .Z(\s9.addr [55]) );
  CAN2XL U6367 ( .A(\s9.addr[7] ), .B(n4164), .Z(\s9.addr [50]) );
  CANR2X1 U6368 ( .A(n3431), .B(\m1.addrM64 [47]), .C(\m3.addrM64 [47]), .D(
        n3289), .Z(n3297) );
  CNR2IX1 U6369 ( .B(\m5.addrM64 [47]), .A(n3432), .Z(n3290) );
  CANR1X1 U6370 ( .A(n3434), .B(\m0.addrM64 [47]), .C(n3290), .Z(n3296) );
  CND2X1 U6371 ( .A(n3435), .B(\m6.addrM64 [47]), .Z(n3292) );
  CND2X1 U6372 ( .A(n3436), .B(\m2.addrM64 [47]), .Z(n3291) );
  CND2X1 U6373 ( .A(n3292), .B(n3291), .Z(n3294) );
  CNR2IX1 U6374 ( .B(\m4.addrM64 [47]), .A(n3439), .Z(n3293) );
  CNR2X1 U6375 ( .A(n3294), .B(n3293), .Z(n3295) );
  CND3X2 U6376 ( .A(n3297), .B(n3296), .C(n3295), .Z(n4146) );
  CAN2XL U6377 ( .A(\s9.addr[16] ), .B(n4146), .Z(\s9.addr [47]) );
  CIVX2 U6378 ( .A(n3470), .Z(n4324) );
  CNR2X1 U6379 ( .A(n3298), .B(n4324), .Z(\s9.addr [44]) );
  CND2XL U6380 ( .A(n3299), .B(\m3.addrM64 [40]), .Z(n3302) );
  CND2X1 U6381 ( .A(n3434), .B(\m0.addrM64 [40]), .Z(n3301) );
  CND2X1 U6382 ( .A(n3431), .B(\m1.addrM64 [40]), .Z(n3300) );
  CAN3X2 U6383 ( .A(n3302), .B(n3301), .C(n3300), .Z(n3310) );
  CIVX2 U6384 ( .A(\m5.addrM64 [40]), .Z(n3304) );
  CND2X1 U6385 ( .A(n3435), .B(\m6.addrM64 [40]), .Z(n3303) );
  CND2X1 U6386 ( .A(n3436), .B(\m2.addrM64 [40]), .Z(n3306) );
  CND2XL U6387 ( .A(n3424), .B(\m4.addrM64 [40]), .Z(n3305) );
  CND2X1 U6388 ( .A(n3306), .B(n3305), .Z(n3307) );
  CNR2X1 U6389 ( .A(n3308), .B(n3307), .Z(n3309) );
  CAN2XL U6390 ( .A(\s9.addr[7] ), .B(n3486), .Z(\s9.addr [40]) );
  CAN2XL U6391 ( .A(\s3.addr[14] ), .B(n4166), .Z(\s3.addr [52]) );
  CAN2XL U6392 ( .A(\s9.addr[8] ), .B(n4171), .Z(\s9.SbusIn [32]) );
  CAN2XL U6393 ( .A(\s9.addr[8] ), .B(n4119), .Z(\s9.SbusIn [31]) );
  CAN2XL U6394 ( .A(\s9.addr[16] ), .B(n4147), .Z(\s9.SbusIn [26]) );
  CAN2XL U6395 ( .A(\s6.addr [17]), .B(n4126), .Z(\s6.SbusIn [62]) );
  CAN2XL U6396 ( .A(\s6.addr [17]), .B(n4170), .Z(\s6.SbusIn [53]) );
  CAN2XL U6397 ( .A(\s9.addr[16] ), .B(n4152), .Z(\s9.SbusIn [19]) );
  CND2X1 U6398 ( .A(n3434), .B(\m0.DoutM [52]), .Z(n3312) );
  CND2XL U6399 ( .A(n3436), .B(\m2.DoutM [52]), .Z(n3311) );
  CND2X1 U6400 ( .A(n3312), .B(n3311), .Z(n3314) );
  CNR2X1 U6401 ( .A(n3314), .B(n3313), .Z(n3318) );
  CANR2X1 U6402 ( .A(n3431), .B(\m1.DoutM [52]), .C(\m3.DoutM [52]), .D(n3420), 
        .Z(n3317) );
  CNR2IX1 U6403 ( .B(\m4.DoutM [52]), .A(n3439), .Z(n3315) );
  CIVX2 U6404 ( .A(n3315), .Z(n3316) );
  CND3X2 U6405 ( .A(n3318), .B(n3317), .C(n3316), .Z(n3466) );
  CAN2XL U6406 ( .A(\s6.addr [17]), .B(n3466), .Z(\s6.SbusIn [52]) );
  CAN2XL U6407 ( .A(\s9.addr[8] ), .B(n3487), .Z(\s9.SbusIn [16]) );
  CAN2XL U6408 ( .A(\s7.en ), .B(n4122), .Z(\s7.addr [43]) );
  CAN2XL U6409 ( .A(n5590), .B(n4154), .Z(\s9.SbusIn [7]) );
  CND2X1 U6410 ( .A(n3420), .B(\m3.DoutM [45]), .Z(n3321) );
  CND2X1 U6411 ( .A(n3434), .B(\m0.DoutM [45]), .Z(n3320) );
  CND2X1 U6412 ( .A(n3431), .B(\m1.DoutM [45]), .Z(n3319) );
  CAN3X2 U6413 ( .A(n3321), .B(n3320), .C(n3319), .Z(n3329) );
  CIVX2 U6414 ( .A(\m5.DoutM [45]), .Z(n3323) );
  CND2X1 U6415 ( .A(n3435), .B(\m6.DoutM [45]), .Z(n3322) );
  CIVX2 U6416 ( .A(\m4.DoutM [45]), .Z(n3325) );
  CND2X1 U6417 ( .A(n3436), .B(\m2.DoutM [45]), .Z(n3324) );
  CNR2X1 U6418 ( .A(n3327), .B(n3326), .Z(n3328) );
  CND2X2 U6419 ( .A(n3329), .B(n3328), .Z(n4129) );
  CAN2XL U6420 ( .A(\s6.addr [17]), .B(n4129), .Z(\s6.SbusIn [45]) );
  CAN2XL U6421 ( .A(\s6.addr [17]), .B(n4146), .Z(\s6.addr [47]) );
  CAN2XL U6422 ( .A(\s6.addr [17]), .B(n4153), .Z(\s6.addr [42]) );
  CAN2XL U6423 ( .A(\s3.addr[14] ), .B(n3456), .Z(\s3.addr [7]) );
  CAN2XL U6424 ( .A(\s6.addr [17]), .B(n3486), .Z(\s6.addr [40]) );
  CAN2XL U6425 ( .A(\s6.addr [17]), .B(n4204), .Z(\s6.addr [38]) );
  CAN2XL U6426 ( .A(\s9.en ), .B(n4129), .Z(\s9.SbusIn [45]) );
  CAN2XL U6427 ( .A(\s6.addr [17]), .B(n3462), .Z(\s6.addr [22]) );
  CAN2XL U6428 ( .A(\s6.addr [17]), .B(n4331), .Z(\s6.addr [20]) );
  CAN2X1 U6429 ( .A(\s3.addr[9] ), .B(n4333), .Z(\s3.addr [3]) );
  CAN2XL U6430 ( .A(\s9.addr[8] ), .B(n4178), .Z(\s9.SbusIn [34]) );
  CIVX4 U6431 ( .A(n3330), .Z(\s13.addr[15] ) );
  CAN2X1 U6432 ( .A(\s13.addr[15] ), .B(n3331), .Z(\s13.SbusIn [38]) );
  CAN2X1 U6433 ( .A(\s13.addr[15] ), .B(n4237), .Z(\s13.SbusIn [35]) );
  CAN2XL U6434 ( .A(\s11.addr[19] ), .B(n4175), .Z(\s11.SbusIn [54]) );
  CIVX12 U6435 ( .A(n3453), .Z(\s1.addr[15] ) );
  CAN2XL U6436 ( .A(\s1.addr[15] ), .B(n4127), .Z(\s1.SbusIn [50]) );
  CAN2XL U6437 ( .A(\s11.addr[19] ), .B(n4126), .Z(\s11.SbusIn [62]) );
  CIVX20 U6438 ( .A(n3417), .Z(n4332) );
  CAN2X1 U6439 ( .A(n4332), .B(n4333), .Z(\s11.addr [3]) );
  CAN2XL U6440 ( .A(\s1.addr[17] ), .B(n3472), .Z(\s1.SbusIn [46]) );
  CAN2X1 U6441 ( .A(\s14.addr[17] ), .B(n4185), .Z(\s14.SbusIn [0]) );
  CAN2XL U6442 ( .A(\s1.addr[17] ), .B(n4331), .Z(\s1.addr [20]) );
  CAN2X1 U6443 ( .A(\s11.addr[19] ), .B(n4195), .Z(\s11.addr [26]) );
  CAN2XL U6444 ( .A(\s1.addr[15] ), .B(n4165), .Z(\s1.addr [51]) );
  CAN2XL U6445 ( .A(\s14.addr[17] ), .B(n4192), .Z(\s14.SbusIn [2]) );
  CAN2XL U6446 ( .A(\s1.addr[15] ), .B(n4149), .Z(\s1.SbusIn [24]) );
  CAN2XL U6447 ( .A(\s1.addr[17] ), .B(n4129), .Z(\s1.SbusIn [45]) );
  CAN2XL U6448 ( .A(\s1.addr[17] ), .B(n4166), .Z(\s1.addr [52]) );
  CAN2X1 U6449 ( .A(\s11.en ), .B(n4339), .Z(\s11.addr [1]) );
  CAN2XL U6450 ( .A(\s1.addr[17] ), .B(n4167), .Z(\s1.SbusIn [60]) );
  CAN2XL U6451 ( .A(\s1.addr[17] ), .B(n4143), .Z(\s1.SbusIn [40]) );
  CAN2XL U6452 ( .A(\s1.addr[15] ), .B(n3464), .Z(\s1.addr [37]) );
  CAN2XL U6453 ( .A(\s1.addr[15] ), .B(n4126), .Z(\s1.SbusIn [62]) );
  CAN2X1 U6454 ( .A(\s1.en ), .B(n4339), .Z(\s1.addr [1]) );
  CAN2X1 U6455 ( .A(\s1.addr [19]), .B(n4333), .Z(\s1.addr [3]) );
  CAN2XL U6456 ( .A(\s1.addr[17] ), .B(n3480), .Z(\s1.SbusIn [49]) );
  CAN2XL U6457 ( .A(\s11.addr[19] ), .B(n4331), .Z(\s11.addr [20]) );
  CAN2X1 U6458 ( .A(n4332), .B(n3455), .Z(\s11.addr [9]) );
  CAN2XL U6459 ( .A(\s14.addr[17] ), .B(n4179), .Z(\s14.addr [33]) );
  CAN2XL U6460 ( .A(\s14.addr[17] ), .B(n4131), .Z(\s14.addr [34]) );
  CAN2XL U6461 ( .A(\s1.addr[15] ), .B(n3473), .Z(\s1.SbusIn [22]) );
  CAN2XL U6462 ( .A(\s1.addr[15] ), .B(n4179), .Z(\s1.addr [33]) );
  CAN2XL U6463 ( .A(\s11.addr[19] ), .B(n4160), .Z(\s11.addr [31]) );
  CND2X1 U6464 ( .A(n3434), .B(\m0.addrM64 [45]), .Z(n3333) );
  CND2XL U6465 ( .A(n3436), .B(\m2.addrM64 [45]), .Z(n3332) );
  CND2X1 U6466 ( .A(n3333), .B(n3332), .Z(n3335) );
  CNR2X1 U6467 ( .A(n3335), .B(n3334), .Z(n3339) );
  CNR2IX1 U6468 ( .B(\m4.addrM64 [45]), .A(n3439), .Z(n3336) );
  CANR1X1 U6469 ( .A(n3431), .B(\m1.addrM64 [45]), .C(n3336), .Z(n3338) );
  CND2X1 U6470 ( .A(n3420), .B(\m3.addrM64 [45]), .Z(n3337) );
  CND3X2 U6471 ( .A(n3339), .B(n3338), .C(n3337), .Z(n4162) );
  CAN2XL U6472 ( .A(\s1.addr[15] ), .B(n4162), .Z(\s1.addr [45]) );
  CAN2XL U6473 ( .A(\s1.addr[17] ), .B(n4150), .Z(\s1.SbusIn [20]) );
  CAN2XL U6474 ( .A(\s14.addr [11]), .B(n4173), .Z(\s14.addr [35]) );
  CAN2XL U6475 ( .A(\s1.addr[17] ), .B(n4122), .Z(\s1.addr [43]) );
  CAN2XL U6476 ( .A(\s11.addr[19] ), .B(n4118), .Z(\s11.addr [23]) );
  CAN2XL U6477 ( .A(\s14.addr[17] ), .B(n3487), .Z(\s14.SbusIn [16]) );
  CAN2XL U6478 ( .A(\s1.addr[15] ), .B(n4117), .Z(\s1.SbusIn [28]) );
  CAN2XL U6479 ( .A(\s1.addr[17] ), .B(n4163), .Z(\s1.SbusIn [51]) );
  CAN2XL U6480 ( .A(\s1.addr[17] ), .B(n4146), .Z(\s1.addr [47]) );
  CAN2XL U6481 ( .A(\s1.addr[15] ), .B(n4197), .Z(\s1.SbusIn [29]) );
  CAN2X1 U6482 ( .A(\s11.addr[19] ), .B(n3456), .Z(\s11.addr [7]) );
  CAN2XL U6483 ( .A(\s1.addr[17] ), .B(n4145), .Z(\s1.SbusIn [30]) );
  CAN2X1 U6484 ( .A(\s1.addr[15] ), .B(n4153), .Z(\s1.addr [42]) );
  CAN2X1 U6485 ( .A(\s1.addr[17] ), .B(n4119), .Z(\s1.SbusIn [31]) );
  CAN2XL U6486 ( .A(\s1.addr[15] ), .B(n3487), .Z(\s1.SbusIn [16]) );
  CND2X1 U6487 ( .A(n3434), .B(\m0.DoutM [56]), .Z(n3341) );
  CND2XL U6488 ( .A(n3436), .B(\m2.DoutM [56]), .Z(n3340) );
  CND2X1 U6489 ( .A(n3341), .B(n3340), .Z(n3345) );
  CIVX2 U6490 ( .A(\m5.DoutM [56]), .Z(n3343) );
  CND2X1 U6491 ( .A(n3435), .B(\m6.DoutM [56]), .Z(n3342) );
  CNR2X1 U6492 ( .A(n3345), .B(n3344), .Z(n3349) );
  CANR2X1 U6493 ( .A(n3431), .B(\m1.DoutM [56]), .C(\m3.DoutM [56]), .D(n3361), 
        .Z(n3348) );
  CNR2IX1 U6494 ( .B(\m4.DoutM [56]), .A(n3439), .Z(n3346) );
  CIVX2 U6495 ( .A(n3346), .Z(n3347) );
  CAN2XL U6496 ( .A(\s11.addr[19] ), .B(n4159), .Z(\s11.SbusIn [56]) );
  CAN2XL U6497 ( .A(\s1.addr[17] ), .B(n3471), .Z(\s1.addr [41]) );
  CAN2XL U6498 ( .A(\s11.addr[19] ), .B(n4199), .Z(\s11.addr [24]) );
  CAN2XL U6499 ( .A(\s1.addr[15] ), .B(n4123), .Z(\s1.SbusIn [13]) );
  CAN2XL U6500 ( .A(\s1.addr[17] ), .B(n4199), .Z(\s1.addr [24]) );
  CAN2X1 U6501 ( .A(\s14.addr [11]), .B(n4339), .Z(\s14.addr [1]) );
  CAN2XL U6502 ( .A(\s1.addr[17] ), .B(n4157), .Z(\s1.addr [32]) );
  CAN2XL U6503 ( .A(\s1.addr[15] ), .B(n3481), .Z(\s1.SbusIn [12]) );
  CAN2XL U6504 ( .A(\s14.addr[17] ), .B(n4154), .Z(\s14.SbusIn [7]) );
  CND2XL U6505 ( .A(n3431), .B(\m1.addrM64 [25]), .Z(n3351) );
  CND2XL U6506 ( .A(n3436), .B(\m2.addrM64 [25]), .Z(n3350) );
  CND2X1 U6507 ( .A(n3351), .B(n3350), .Z(n3353) );
  CNR2IX1 U6508 ( .B(\m4.addrM64 [25]), .A(n3439), .Z(n3352) );
  CNR2X1 U6509 ( .A(n3353), .B(n3352), .Z(n3357) );
  CANR2X1 U6510 ( .A(n3420), .B(\m3.addrM64 [25]), .C(\m6.addrM64 [25]), .D(
        n3435), .Z(n3356) );
  CNR2IX1 U6511 ( .B(\m5.addrM64 [25]), .A(n3432), .Z(n3354) );
  CANR1X1 U6512 ( .A(n3434), .B(\m0.addrM64 [25]), .C(n3354), .Z(n3355) );
  CND3X2 U6513 ( .A(n3357), .B(n3356), .C(n3355), .Z(n4328) );
  CAN2XL U6514 ( .A(\s11.addr[19] ), .B(n4328), .Z(\s11.addr [25]) );
  CAN2XL U6515 ( .A(\s1.addr[17] ), .B(n4215), .Z(\s1.SbusIn [36]) );
  CAN2XL U6516 ( .A(\s1.addr[17] ), .B(n3462), .Z(\s1.addr [22]) );
  CAN2XL U6517 ( .A(\s14.addr[17] ), .B(n4200), .Z(\s14.SbusIn [3]) );
  CAN2XL U6518 ( .A(n4050), .B(n3482), .Z(\s10.addr [60]) );
  CAN2XL U6519 ( .A(n4050), .B(n4197), .Z(\s10.SbusIn [29]) );
  CAN2XL U6520 ( .A(n4050), .B(n4145), .Z(\s10.SbusIn [30]) );
  CAN2XL U6521 ( .A(\s11.en ), .B(n4190), .Z(\s11.SbusIn [1]) );
  CAN2XL U6522 ( .A(\s11.en ), .B(n4169), .Z(\s11.SbusIn [15]) );
  CAN2XL U6523 ( .A(n4050), .B(n4115), .Z(\s10.SbusIn [10]) );
  CAN2XL U6524 ( .A(\s10.addr[9] ), .B(n4172), .Z(\s10.SbusIn [17]) );
  CAN2XL U6525 ( .A(\s10.addr[9] ), .B(n4193), .Z(\s10.SbusIn [9]) );
  CAN2XL U6526 ( .A(\s10.addr[9] ), .B(n4116), .Z(\s10.SbusIn [8]) );
  CAN2XL U6527 ( .A(n4050), .B(n4154), .Z(\s10.SbusIn [7]) );
  CAN2XL U6528 ( .A(\s11.en ), .B(n4200), .Z(\s11.SbusIn [3]) );
  CAN2XL U6529 ( .A(\s10.addr[9] ), .B(n4243), .Z(\s10.SbusIn [4]) );
  CAN2XL U6530 ( .A(\s10.addr[9] ), .B(n4175), .Z(\s10.SbusIn [54]) );
  CAN2XL U6531 ( .A(\s9.addr[16] ), .B(n4169), .Z(\s9.SbusIn [15]) );
  CNR2IX1 U6532 ( .B(\m5.DoutM [57]), .A(n3432), .Z(n3358) );
  CNR2IX1 U6533 ( .B(\m4.DoutM [57]), .A(n3439), .Z(n3359) );
  CIVX2 U6534 ( .A(n3359), .Z(n3364) );
  CAN2X1 U6535 ( .A(n3435), .B(\m6.DoutM [57]), .Z(n3360) );
  CANR2X1 U6536 ( .A(n3434), .B(\m0.DoutM [57]), .C(n3436), .D(\m2.DoutM [57]), 
        .Z(n3362) );
  CND4X2 U6537 ( .A(n3365), .B(n3364), .C(n3363), .D(n3362), .Z(n4161) );
  CAN2XL U6538 ( .A(n4050), .B(n4161), .Z(\s10.SbusIn [57]) );
  CAN2XL U6539 ( .A(n4050), .B(n4168), .Z(\s10.SbusIn [58]) );
  CAN2XL U6540 ( .A(\s11.addr[19] ), .B(n3460), .Z(\s11.SbusIn [27]) );
  CAN2XL U6541 ( .A(\s11.en ), .B(n4117), .Z(\s11.SbusIn [28]) );
  CAN2XL U6542 ( .A(\s11.addr[19] ), .B(n4143), .Z(\s11.SbusIn [40]) );
  CAN2XL U6543 ( .A(\s9.addr[7] ), .B(n4143), .Z(\s9.SbusIn [40]) );
  CAN2XL U6544 ( .A(\s9.addr[8] ), .B(n4132), .Z(\s9.SbusIn [43]) );
  CAN2XL U6545 ( .A(\s11.addr[19] ), .B(n4197), .Z(\s11.SbusIn [29]) );
  CAN2XL U6546 ( .A(\s11.en ), .B(n3469), .Z(\s11.SbusIn [5]) );
  CAN2XL U6547 ( .A(\s9.addr[16] ), .B(n4161), .Z(\s9.SbusIn [57]) );
  CAN2XL U6548 ( .A(n4050), .B(n4125), .Z(\s10.SbusIn [61]) );
  CAN2XL U6549 ( .A(\s11.addr[19] ), .B(n4119), .Z(\s11.SbusIn [31]) );
  CAN2XL U6550 ( .A(\s9.addr[16] ), .B(n4167), .Z(\s9.SbusIn [60]) );
  CAN2X1 U6551 ( .A(\s9.addr [15]), .B(n4334), .Z(\s9.addr [4]) );
  CAN2XL U6552 ( .A(\s11.addr[19] ), .B(n4329), .Z(\s11.SbusIn [6]) );
  CAN2XL U6553 ( .A(\s11.addr[19] ), .B(n4196), .Z(\s11.SbusIn [37]) );
  CAN2XL U6554 ( .A(\s9.addr[16] ), .B(n4155), .Z(\s9.addr [49]) );
  CAN2XL U6555 ( .A(n5590), .B(n4137), .Z(\s9.addr [48]) );
  CAN2XL U6556 ( .A(\s10.addr[9] ), .B(n4123), .Z(\s10.SbusIn [13]) );
  CAN2XL U6557 ( .A(\s1.addr[17] ), .B(n4151), .Z(\s1.addr [61]) );
  CAN2XL U6558 ( .A(\s11.addr[19] ), .B(n4129), .Z(\s11.SbusIn [45]) );
  CAN2XL U6559 ( .A(\s11.en ), .B(n4138), .Z(\s11.SbusIn [44]) );
  CAN2XL U6560 ( .A(\s1.addr[15] ), .B(n3482), .Z(\s1.addr [60]) );
  CAN2XL U6561 ( .A(\s1.addr[15] ), .B(n4193), .Z(\s1.SbusIn [9]) );
  CAN2XL U6562 ( .A(n4050), .B(n4141), .Z(\s10.SbusIn [25]) );
  CAN2XL U6563 ( .A(n4050), .B(n4173), .Z(\s10.addr [35]) );
  CAN2XL U6564 ( .A(\s1.addr[17] ), .B(n4242), .Z(\s1.addr [56]) );
  CAN2XL U6565 ( .A(\s1.addr[17] ), .B(n3477), .Z(\s1.addr [59]) );
  CAN2XL U6566 ( .A(\s11.addr[19] ), .B(n4180), .Z(\s11.SbusIn [18]) );
  CAN2XL U6567 ( .A(n4050), .B(n3464), .Z(\s10.addr [37]) );
  CND2X1 U6568 ( .A(n3434), .B(\m0.DoutM [47]), .Z(n3367) );
  CND2XL U6569 ( .A(n3436), .B(\m2.DoutM [47]), .Z(n3366) );
  CND2X1 U6570 ( .A(n3367), .B(n3366), .Z(n3369) );
  CNR2X1 U6571 ( .A(n3369), .B(n3368), .Z(n3374) );
  CNR2IX1 U6572 ( .B(\m4.DoutM [47]), .A(n3439), .Z(n3370) );
  CANR1X1 U6573 ( .A(n3431), .B(\m1.DoutM [47]), .C(n3370), .Z(n3373) );
  CND2X2 U6574 ( .A(n3371), .B(\m3.DoutM [47]), .Z(n3372) );
  CND3X2 U6575 ( .A(n3374), .B(n3373), .C(n3372), .Z(n4139) );
  CAN2XL U6576 ( .A(\s11.addr[19] ), .B(n4139), .Z(\s11.SbusIn [47]) );
  CNR2IX1 U6577 ( .B(n4196), .A(n3375), .Z(\s13.SbusIn [37]) );
  CAN2XL U6578 ( .A(\s10.addr[9] ), .B(n4150), .Z(\s10.SbusIn [20]) );
  CAN2XL U6579 ( .A(n4050), .B(n4124), .Z(\s10.addr [36]) );
  CNR2IX1 U6580 ( .B(n3376), .A(n3375), .Z(\s13.SbusIn [36]) );
  CAN2XL U6581 ( .A(\s1.addr[17] ), .B(n4201), .Z(\s1.addr [55]) );
  CAN2XL U6582 ( .A(\s11.addr[19] ), .B(n4172), .Z(\s11.SbusIn [17]) );
  CAN2X1 U6583 ( .A(n4050), .B(n4177), .Z(\s10.addr [39]) );
  CIVX12 U6584 ( .A(n3449), .Z(\s3.addr [18]) );
  CNR2X1 U6585 ( .A(n3446), .B(n4326), .Z(\s1.addr [6]) );
  CIVX8 U6586 ( .A(n3377), .Z(\s2.addr[19] ) );
  CNR2IX1 U6587 ( .B(n3462), .A(n3378), .Z(\s10.addr [22]) );
  CNR2XL U6588 ( .A(n3379), .B(n5580), .Z(\m3.MinData [56]) );
  CNR2XL U6589 ( .A(n3379), .B(n5581), .Z(\m3.MinData [57]) );
  CNR2XL U6590 ( .A(n3379), .B(n5587), .Z(\m3.MinData [63]) );
  CNR2XL U6591 ( .A(n3379), .B(n5582), .Z(\m3.MinData [58]) );
  CNR2XL U6592 ( .A(n3379), .B(n5586), .Z(\m3.MinData [62]) );
  CNR2XL U6593 ( .A(n3379), .B(n5583), .Z(\m3.MinData [59]) );
  CNR2XL U6594 ( .A(n3379), .B(n5584), .Z(\m3.MinData [60]) );
  CNR2XL U6595 ( .A(n3379), .B(n5585), .Z(\m3.MinData [61]) );
  CNR2XL U6596 ( .A(n3379), .B(n5579), .Z(\m3.MinData [55]) );
  CNR2XL U6597 ( .A(n3379), .B(n5567), .Z(\m3.MinData [44]) );
  CNR2XL U6598 ( .A(n3379), .B(n5578), .Z(\m3.MinData [54]) );
  CNR2XL U6599 ( .A(n3379), .B(n5577), .Z(\m3.MinData [53]) );
  CNR2XL U6600 ( .A(n3379), .B(n5568), .Z(\m3.MinData [45]) );
  CNR2XL U6601 ( .A(n3379), .B(n5569), .Z(\m3.MinData [46]) );
  CNR2XL U6602 ( .A(n3379), .B(n5576), .Z(\m3.MinData [52]) );
  CNR2XL U6603 ( .A(n3379), .B(n5570), .Z(\m3.MinData [47]) );
  CNR2XL U6604 ( .A(n3379), .B(n5571), .Z(\m3.MinData [48]) );
  CNR2XL U6605 ( .A(n3379), .B(n5575), .Z(\m3.MinData [51]) );
  CNR2XL U6606 ( .A(n3379), .B(n5572), .Z(\m3.MinData [49]) );
  CNR2XL U6607 ( .A(n3379), .B(n5574), .Z(\m3.MinData [50]) );
  CNR2XL U6608 ( .A(n3379), .B(n5530), .Z(\m3.MinData [7]) );
  CNR2XL U6609 ( .A(n3379), .B(n5552), .Z(\m3.MinData [29]) );
  CNR2XL U6610 ( .A(n3379), .B(n5531), .Z(\m3.MinData [8]) );
  CNR2XL U6611 ( .A(n3379), .B(n5551), .Z(\m3.MinData [28]) );
  CNR2XL U6612 ( .A(n3379), .B(n5532), .Z(\m3.MinData [9]) );
  CNR2XL U6613 ( .A(n3379), .B(n5550), .Z(\m3.MinData [27]) );
  CNR2XL U6614 ( .A(n3379), .B(n5549), .Z(\m3.MinData [26]) );
  CNR2XL U6615 ( .A(n3379), .B(n5533), .Z(\m3.MinData [10]) );
  CNR2XL U6616 ( .A(n3379), .B(n5548), .Z(\m3.MinData [25]) );
  CNR2XL U6617 ( .A(n3379), .B(n5547), .Z(\m3.MinData [24]) );
  CNR2XL U6618 ( .A(n3379), .B(n5546), .Z(\m3.MinData [23]) );
  CNR2XL U6619 ( .A(n3379), .B(n5534), .Z(\m3.MinData [11]) );
  CNR2XL U6620 ( .A(n3379), .B(n5545), .Z(\m3.MinData [22]) );
  CNR2XL U6621 ( .A(n3379), .B(n5535), .Z(\m3.MinData [12]) );
  CNR2XL U6622 ( .A(n3379), .B(n5544), .Z(\m3.MinData [21]) );
  CNR2XL U6623 ( .A(n3379), .B(n5543), .Z(\m3.MinData [20]) );
  CNR2XL U6624 ( .A(n3379), .B(n5542), .Z(\m3.MinData [19]) );
  CNR2XL U6625 ( .A(n3379), .B(n5541), .Z(\m3.MinData [18]) );
  CNR2XL U6626 ( .A(n3379), .B(n5540), .Z(\m3.MinData [17]) );
  CNR2XL U6627 ( .A(n3379), .B(n5539), .Z(\m3.MinData [16]) );
  CNR2XL U6628 ( .A(n3379), .B(n5536), .Z(\m3.MinData [13]) );
  CNR2XL U6629 ( .A(n3379), .B(n5538), .Z(\m3.MinData [15]) );
  CNR2XL U6630 ( .A(n3379), .B(n5537), .Z(\m3.MinData [14]) );
  CNR2XL U6631 ( .A(n3379), .B(n5566), .Z(\m3.MinData [43]) );
  CNR2XL U6632 ( .A(n3379), .B(n5565), .Z(\m3.MinData [42]) );
  CNR2XL U6633 ( .A(n3379), .B(n5564), .Z(\m3.MinData [41]) );
  CNR2XL U6634 ( .A(n3379), .B(n5563), .Z(\m3.MinData [40]) );
  CNR2XL U6635 ( .A(n3379), .B(n5562), .Z(\m3.MinData [39]) );
  CNR2XL U6636 ( .A(n3379), .B(n5561), .Z(\m3.MinData [38]) );
  CNR2XL U6637 ( .A(n3379), .B(n5560), .Z(\m3.MinData [37]) );
  CNR2XL U6638 ( .A(n3379), .B(n5525), .Z(\m3.MinData [2]) );
  CNR2XL U6639 ( .A(n3379), .B(n5526), .Z(\m3.MinData [3]) );
  CNR2XL U6640 ( .A(n3379), .B(n5559), .Z(\m3.MinData [36]) );
  CNR2XL U6641 ( .A(n3379), .B(n5558), .Z(\m3.MinData [35]) );
  CNR2XL U6642 ( .A(n3379), .B(n5528), .Z(\m3.MinData [5]) );
  CNR2XL U6643 ( .A(n3379), .B(n5557), .Z(\m3.MinData [34]) );
  CNR2XL U6644 ( .A(n3379), .B(n5556), .Z(\m3.MinData [33]) );
  CNR2XL U6645 ( .A(n3379), .B(n5527), .Z(\m3.MinData [4]) );
  CNR2XL U6646 ( .A(n3379), .B(n5553), .Z(\m3.MinData [30]) );
  CNR2XL U6647 ( .A(n3379), .B(n5555), .Z(\m3.MinData [32]) );
  CNR2XL U6648 ( .A(n3379), .B(n5523), .Z(\m3.MinData [0]) );
  CNR2XL U6649 ( .A(n3379), .B(n5524), .Z(\m3.MinData [1]) );
  CNR2XL U6650 ( .A(n3379), .B(n5554), .Z(\m3.MinData [31]) );
  CNR2XL U6651 ( .A(n3379), .B(n5529), .Z(\m3.MinData [6]) );
  CNR2XL U6652 ( .A(n3380), .B(n5577), .Z(\m0.MinData [53]) );
  CNR2XL U6653 ( .A(n3380), .B(n5579), .Z(\m0.MinData [55]) );
  CNR2XL U6654 ( .A(n3380), .B(n5576), .Z(\m0.MinData [52]) );
  CNR2XL U6655 ( .A(n3380), .B(n5523), .Z(\m0.MinData [0]) );
  CNR2XL U6656 ( .A(n3380), .B(n5524), .Z(\m0.MinData [1]) );
  CNR2XL U6657 ( .A(n3380), .B(n5525), .Z(\m0.MinData [2]) );
  CNR2XL U6658 ( .A(n3380), .B(n5526), .Z(\m0.MinData [3]) );
  CNR2XL U6659 ( .A(n3380), .B(n5578), .Z(\m0.MinData [54]) );
  CNR2XL U6660 ( .A(n3380), .B(n5527), .Z(\m0.MinData [4]) );
  CNR2XL U6661 ( .A(n3380), .B(n5575), .Z(\m0.MinData [51]) );
  CNR2XL U6662 ( .A(n3380), .B(n5580), .Z(\m0.MinData [56]) );
  CNR2XL U6663 ( .A(n3380), .B(n5581), .Z(\m0.MinData [57]) );
  CNR2XL U6664 ( .A(n3380), .B(n5582), .Z(\m0.MinData [58]) );
  CNR2XL U6665 ( .A(n3380), .B(n5583), .Z(\m0.MinData [59]) );
  CNR2XL U6666 ( .A(n3380), .B(n5559), .Z(\m0.MinData [36]) );
  CNR2XL U6667 ( .A(n3380), .B(n5535), .Z(\m0.MinData [12]) );
  CNR2XL U6668 ( .A(n3380), .B(n5558), .Z(\m0.MinData [35]) );
  CNR2XL U6669 ( .A(n3380), .B(n5534), .Z(\m0.MinData [11]) );
  CNR2XL U6670 ( .A(n3380), .B(n5561), .Z(\m0.MinData [38]) );
  CNR2XL U6671 ( .A(n3380), .B(n5557), .Z(\m0.MinData [34]) );
  CNR2XL U6672 ( .A(n3380), .B(n5533), .Z(\m0.MinData [10]) );
  CNR2XL U6673 ( .A(n3380), .B(n5532), .Z(\m0.MinData [9]) );
  CNR2XL U6674 ( .A(n3380), .B(n5556), .Z(\m0.MinData [33]) );
  CNR2XL U6675 ( .A(n3380), .B(n5562), .Z(\m0.MinData [39]) );
  CNR2XL U6676 ( .A(n3380), .B(n5531), .Z(\m0.MinData [8]) );
  CNR2XL U6677 ( .A(n3380), .B(n5555), .Z(\m0.MinData [32]) );
  CNR2XL U6678 ( .A(n3380), .B(n5563), .Z(\m0.MinData [40]) );
  CNR2XL U6679 ( .A(n3380), .B(n5530), .Z(\m0.MinData [7]) );
  CNR2XL U6680 ( .A(n3380), .B(n5554), .Z(\m0.MinData [31]) );
  CNR2XL U6681 ( .A(n3380), .B(n5564), .Z(\m0.MinData [41]) );
  CNR2XL U6682 ( .A(n3380), .B(n5529), .Z(\m0.MinData [6]) );
  CNR2XL U6683 ( .A(n3380), .B(n5565), .Z(\m0.MinData [42]) );
  CNR2XL U6684 ( .A(n3380), .B(n5542), .Z(\m0.MinData [19]) );
  CNR2XL U6685 ( .A(n3380), .B(n5528), .Z(\m0.MinData [5]) );
  CNR2XL U6686 ( .A(n3380), .B(n5543), .Z(\m0.MinData [20]) );
  CNR2XL U6687 ( .A(n3380), .B(n5544), .Z(\m0.MinData [21]) );
  CNR2XL U6688 ( .A(n3380), .B(n5545), .Z(\m0.MinData [22]) );
  CNR2XL U6689 ( .A(n3380), .B(n5546), .Z(\m0.MinData [23]) );
  CNR2XL U6690 ( .A(n3380), .B(n5567), .Z(\m0.MinData [44]) );
  CNR2XL U6691 ( .A(n3380), .B(n5536), .Z(\m0.MinData [13]) );
  CNR2XL U6692 ( .A(n3380), .B(n5560), .Z(\m0.MinData [37]) );
  CNR2XL U6693 ( .A(n3380), .B(n5537), .Z(\m0.MinData [14]) );
  CNR2XL U6694 ( .A(n3380), .B(n5547), .Z(\m0.MinData [24]) );
  CNR2XL U6695 ( .A(n3380), .B(n5574), .Z(\m0.MinData [50]) );
  CNR2XL U6696 ( .A(n3380), .B(n5548), .Z(\m0.MinData [25]) );
  CNR2XL U6697 ( .A(n3380), .B(n5552), .Z(\m0.MinData [29]) );
  CNR2XL U6698 ( .A(n3380), .B(n5549), .Z(\m0.MinData [26]) );
  CNR2XL U6699 ( .A(n3380), .B(n5566), .Z(\m0.MinData [43]) );
  CNR2XL U6700 ( .A(n3380), .B(n5553), .Z(\m0.MinData [30]) );
  CNR2XL U6701 ( .A(n3380), .B(n5539), .Z(\m0.MinData [16]) );
  CNR2XL U6702 ( .A(n3380), .B(n5538), .Z(\m0.MinData [15]) );
  CNR2XL U6703 ( .A(n3380), .B(n5550), .Z(\m0.MinData [27]) );
  CNR2XL U6704 ( .A(n3380), .B(n5540), .Z(\m0.MinData [17]) );
  CNR2XL U6705 ( .A(n3380), .B(n5551), .Z(\m0.MinData [28]) );
  CNR2XL U6706 ( .A(n3380), .B(n5541), .Z(\m0.MinData [18]) );
  CNR2XL U6707 ( .A(n3381), .B(n5554), .Z(\m6.MinData [31]) );
  CNR2XL U6708 ( .A(n3381), .B(n5557), .Z(\m6.MinData [34]) );
  CNR2XL U6709 ( .A(n3381), .B(n5553), .Z(\m6.MinData [30]) );
  CNR2XL U6710 ( .A(n3381), .B(n5552), .Z(\m6.MinData [29]) );
  CNR2XL U6711 ( .A(n3381), .B(n5555), .Z(\m6.MinData [32]) );
  CNR2XL U6712 ( .A(n3381), .B(n5556), .Z(\m6.MinData [33]) );
  CNR2XL U6713 ( .A(n3381), .B(n5551), .Z(\m6.MinData [28]) );
  CNR2XL U6714 ( .A(n3381), .B(n5550), .Z(\m6.MinData [27]) );
  CNR2XL U6715 ( .A(n3381), .B(n5549), .Z(\m6.MinData [26]) );
  CNR2XL U6716 ( .A(n3381), .B(n5548), .Z(\m6.MinData [25]) );
  CNR2XL U6717 ( .A(n3381), .B(n5547), .Z(\m6.MinData [24]) );
  CNR2XL U6718 ( .A(n3381), .B(n5546), .Z(\m6.MinData [23]) );
  CNR2XL U6719 ( .A(n3381), .B(n5545), .Z(\m6.MinData [22]) );
  CNR2XL U6720 ( .A(n3381), .B(n5544), .Z(\m6.MinData [21]) );
  CNR2XL U6721 ( .A(n3381), .B(n5543), .Z(\m6.MinData [20]) );
  CNR2XL U6722 ( .A(n3381), .B(n5542), .Z(\m6.MinData [19]) );
  CNR2XL U6723 ( .A(n3381), .B(n5541), .Z(\m6.MinData [18]) );
  CNR2XL U6724 ( .A(n3381), .B(n5540), .Z(\m6.MinData [17]) );
  CNR2XL U6725 ( .A(n3381), .B(n5539), .Z(\m6.MinData [16]) );
  CNR2XL U6726 ( .A(n3381), .B(n5538), .Z(\m6.MinData [15]) );
  CNR2XL U6727 ( .A(n3381), .B(n5537), .Z(\m6.MinData [14]) );
  CNR2XL U6728 ( .A(n3381), .B(n5536), .Z(\m6.MinData [13]) );
  CNR2XL U6729 ( .A(n3381), .B(n5535), .Z(\m6.MinData [12]) );
  CNR2XL U6730 ( .A(n3381), .B(n5581), .Z(\m6.MinData [57]) );
  CNR2XL U6731 ( .A(n3381), .B(n5583), .Z(\m6.MinData [59]) );
  CNR2XL U6732 ( .A(n3381), .B(n5580), .Z(\m6.MinData [56]) );
  CNR2XL U6733 ( .A(n3381), .B(n5579), .Z(\m6.MinData [55]) );
  CNR2XL U6734 ( .A(n3381), .B(n5578), .Z(\m6.MinData [54]) );
  CNR2XL U6735 ( .A(n3381), .B(n5577), .Z(\m6.MinData [53]) );
  CNR2XL U6736 ( .A(n3381), .B(n5576), .Z(\m6.MinData [52]) );
  CNR2XL U6737 ( .A(n3381), .B(n5575), .Z(\m6.MinData [51]) );
  CNR2XL U6738 ( .A(n3381), .B(n5574), .Z(\m6.MinData [50]) );
  CNR2XL U6739 ( .A(n3381), .B(n5567), .Z(\m6.MinData [44]) );
  CNR2XL U6740 ( .A(n3381), .B(n5566), .Z(\m6.MinData [43]) );
  CNR2XL U6741 ( .A(n3381), .B(n5565), .Z(\m6.MinData [42]) );
  CNR2XL U6742 ( .A(n3381), .B(n5582), .Z(\m6.MinData [58]) );
  CNR2XL U6743 ( .A(n3381), .B(n5564), .Z(\m6.MinData [41]) );
  CNR2XL U6744 ( .A(n3381), .B(n5563), .Z(\m6.MinData [40]) );
  CNR2XL U6745 ( .A(n3381), .B(n5562), .Z(\m6.MinData [39]) );
  CNR2XL U6746 ( .A(n3381), .B(n5561), .Z(\m6.MinData [38]) );
  CNR2XL U6747 ( .A(n3381), .B(n5560), .Z(\m6.MinData [37]) );
  CNR2XL U6748 ( .A(n3381), .B(n5559), .Z(\m6.MinData [36]) );
  CNR2XL U6749 ( .A(n3381), .B(n5558), .Z(\m6.MinData [35]) );
  CNR2XL U6750 ( .A(n3381), .B(n5532), .Z(\m6.MinData [9]) );
  CNR2XL U6751 ( .A(n3381), .B(n5531), .Z(\m6.MinData [8]) );
  CNR2XL U6752 ( .A(n3381), .B(n5530), .Z(\m6.MinData [7]) );
  CNR2XL U6753 ( .A(n3381), .B(n5529), .Z(\m6.MinData [6]) );
  CNR2XL U6754 ( .A(n3381), .B(n5528), .Z(\m6.MinData [5]) );
  CNR2XL U6755 ( .A(n3381), .B(n5527), .Z(\m6.MinData [4]) );
  CNR2XL U6756 ( .A(n3381), .B(n5526), .Z(\m6.MinData [3]) );
  CNR2XL U6757 ( .A(n3381), .B(n5525), .Z(\m6.MinData [2]) );
  CNR2XL U6758 ( .A(n3381), .B(n5524), .Z(\m6.MinData [1]) );
  CNR2XL U6759 ( .A(n3381), .B(n5523), .Z(\m6.MinData [0]) );
  CNR2XL U6760 ( .A(n3381), .B(n5534), .Z(\m6.MinData [11]) );
  CNR2XL U6761 ( .A(n3381), .B(n5533), .Z(\m6.MinData [10]) );
  CNR2XL U6762 ( .A(n3382), .B(n5558), .Z(\m2.MinData [35]) );
  CNR2XL U6763 ( .A(n3382), .B(n5557), .Z(\m2.MinData [34]) );
  CNR2XL U6764 ( .A(n3382), .B(n5556), .Z(\m2.MinData [33]) );
  CNR2XL U6765 ( .A(n3382), .B(n5559), .Z(\m2.MinData [36]) );
  CNR2XL U6766 ( .A(n3382), .B(n5555), .Z(\m2.MinData [32]) );
  CNR2XL U6767 ( .A(n3382), .B(n5554), .Z(\m2.MinData [31]) );
  CNR2XL U6768 ( .A(n3382), .B(n5553), .Z(\m2.MinData [30]) );
  CNR2XL U6769 ( .A(n3382), .B(n5560), .Z(\m2.MinData [37]) );
  CNR2XL U6770 ( .A(n3382), .B(n5552), .Z(\m2.MinData [29]) );
  CNR2XL U6771 ( .A(n3382), .B(n5551), .Z(\m2.MinData [28]) );
  CNR2XL U6772 ( .A(n3382), .B(n5550), .Z(\m2.MinData [27]) );
  CNR2XL U6773 ( .A(n3382), .B(n5561), .Z(\m2.MinData [38]) );
  CNR2XL U6774 ( .A(n3382), .B(n5549), .Z(\m2.MinData [26]) );
  CNR2XL U6775 ( .A(n3382), .B(n5548), .Z(\m2.MinData [25]) );
  CNR2XL U6776 ( .A(n3382), .B(n5547), .Z(\m2.MinData [24]) );
  CNR2XL U6777 ( .A(n3382), .B(n5546), .Z(\m2.MinData [23]) );
  CNR2XL U6778 ( .A(n3382), .B(n5545), .Z(\m2.MinData [22]) );
  CNR2XL U6779 ( .A(n3382), .B(n5562), .Z(\m2.MinData [39]) );
  CNR2XL U6780 ( .A(n3382), .B(n5544), .Z(\m2.MinData [21]) );
  CNR2XL U6781 ( .A(n3382), .B(n5543), .Z(\m2.MinData [20]) );
  CNR2XL U6782 ( .A(n3382), .B(n5542), .Z(\m2.MinData [19]) );
  CNR2XL U6783 ( .A(n3382), .B(n5541), .Z(\m2.MinData [18]) );
  CNR2XL U6784 ( .A(n3382), .B(n5563), .Z(\m2.MinData [40]) );
  CNR2XL U6785 ( .A(n3382), .B(n5539), .Z(\m2.MinData [16]) );
  CNR2XL U6786 ( .A(n3382), .B(n5564), .Z(\m2.MinData [41]) );
  CNR2XL U6787 ( .A(n3382), .B(n5538), .Z(\m2.MinData [15]) );
  CNR2XL U6788 ( .A(n3382), .B(n5537), .Z(\m2.MinData [14]) );
  CNR2XL U6789 ( .A(n3382), .B(n5536), .Z(\m2.MinData [13]) );
  CNR2XL U6790 ( .A(n3382), .B(n5535), .Z(\m2.MinData [12]) );
  CNR2XL U6791 ( .A(n3382), .B(n5565), .Z(\m2.MinData [42]) );
  CNR2XL U6792 ( .A(n3382), .B(n5534), .Z(\m2.MinData [11]) );
  CNR2XL U6793 ( .A(n3382), .B(n5533), .Z(\m2.MinData [10]) );
  CNR2XL U6794 ( .A(n3382), .B(n5532), .Z(\m2.MinData [9]) );
  CNR2XL U6795 ( .A(n3382), .B(n5531), .Z(\m2.MinData [8]) );
  CNR2XL U6796 ( .A(n3382), .B(n5530), .Z(\m2.MinData [7]) );
  CNR2XL U6797 ( .A(n3382), .B(n5566), .Z(\m2.MinData [43]) );
  CNR2XL U6798 ( .A(n3382), .B(n5567), .Z(\m2.MinData [44]) );
  CNR2XL U6799 ( .A(n3382), .B(n5529), .Z(\m2.MinData [6]) );
  CNR2XL U6800 ( .A(n3382), .B(n5568), .Z(\m2.MinData [45]) );
  CNR2XL U6801 ( .A(n3382), .B(n5528), .Z(\m2.MinData [5]) );
  CNR2XL U6802 ( .A(n3382), .B(n5569), .Z(\m2.MinData [46]) );
  CNR2XL U6803 ( .A(n3382), .B(n5527), .Z(\m2.MinData [4]) );
  CNR2XL U6804 ( .A(n3382), .B(n5526), .Z(\m2.MinData [3]) );
  CNR2XL U6805 ( .A(n3382), .B(n5570), .Z(\m2.MinData [47]) );
  CNR2XL U6806 ( .A(n3382), .B(n5525), .Z(\m2.MinData [2]) );
  CNR2XL U6807 ( .A(n3382), .B(n5571), .Z(\m2.MinData [48]) );
  CNR2XL U6808 ( .A(n3382), .B(n5524), .Z(\m2.MinData [1]) );
  CNR2XL U6809 ( .A(n3382), .B(n5523), .Z(\m2.MinData [0]) );
  CNR2XL U6810 ( .A(n3382), .B(n5572), .Z(\m2.MinData [49]) );
  CNR2XL U6811 ( .A(n3382), .B(n5579), .Z(\m2.MinData [55]) );
  CNR2XL U6812 ( .A(n3382), .B(n5580), .Z(\m2.MinData [56]) );
  CNR2XL U6813 ( .A(n3382), .B(n5581), .Z(\m2.MinData [57]) );
  CNR2XL U6814 ( .A(n3382), .B(n5582), .Z(\m2.MinData [58]) );
  CNR2XL U6815 ( .A(n3382), .B(n5583), .Z(\m2.MinData [59]) );
  CNR2XL U6816 ( .A(n3382), .B(n5540), .Z(\m2.MinData [17]) );
  CNR2XL U6817 ( .A(n3383), .B(n5557), .Z(\m1.MinData [34]) );
  CNR2XL U6818 ( .A(n3383), .B(n5575), .Z(\m1.MinData [51]) );
  CNR2XL U6819 ( .A(n3383), .B(n5559), .Z(\m1.MinData [36]) );
  CNR2XL U6820 ( .A(n3383), .B(n5562), .Z(\m1.MinData [39]) );
  CNR2XL U6821 ( .A(n3383), .B(n5554), .Z(\m1.MinData [31]) );
  CNR2XL U6822 ( .A(n3383), .B(n5563), .Z(\m1.MinData [40]) );
  CNR2XL U6823 ( .A(n3383), .B(n5570), .Z(\m1.MinData [47]) );
  CNR2XL U6824 ( .A(n3383), .B(n5566), .Z(\m1.MinData [43]) );
  CNR2XL U6825 ( .A(n3383), .B(n5530), .Z(\m1.MinData [7]) );
  CNR2XL U6826 ( .A(n3383), .B(n5587), .Z(\m1.MinData [63]) );
  CNR2XL U6827 ( .A(n3383), .B(n5527), .Z(\m1.MinData [4]) );
  CNR2XL U6828 ( .A(n3383), .B(n5526), .Z(\m1.MinData [3]) );
  CNR2XL U6829 ( .A(n3383), .B(n5525), .Z(\m1.MinData [2]) );
  CNR2XL U6830 ( .A(n3383), .B(n5524), .Z(\m1.MinData [1]) );
  CNR2XL U6831 ( .A(n3383), .B(n5584), .Z(\m1.MinData [60]) );
  CNR2XL U6832 ( .A(n3383), .B(n5523), .Z(\m1.MinData [0]) );
  CNR2XL U6833 ( .A(n3383), .B(n5582), .Z(\m1.MinData [58]) );
  CNR2XL U6834 ( .A(n3383), .B(n5545), .Z(\m1.MinData [22]) );
  CNR2XL U6835 ( .A(n3383), .B(n5548), .Z(\m1.MinData [25]) );
  CNR2XL U6836 ( .A(n3383), .B(n5579), .Z(\m1.MinData [55]) );
  CNR2XL U6837 ( .A(n3383), .B(n5578), .Z(\m1.MinData [54]) );
  CNR2XL U6838 ( .A(n3383), .B(n5551), .Z(\m1.MinData [28]) );
  CIVXL U6839 ( .A(n3384), .Z(n3402) );
  CIVX1 U6840 ( .A(\m1.need ), .Z(n3386) );
  CANR3X1 U6841 ( .A(\m2.need ), .B(n3386), .C(\m6.need ), .D(\m0.need ), .Z(
        n3387) );
  CNR2X1 U6842 ( .A(\m3.need ), .B(n3387), .Z(n3388) );
  CNR2X1 U6843 ( .A(n3388), .B(\m4.need ), .Z(n3390) );
  CIVXL U6844 ( .A(n3389), .Z(n3401) );
  COND11X1 U6845 ( .A(n3402), .B(n1846), .C(n3390), .D(n3389), .Z(n3391) );
  CIVX1 U6846 ( .A(n3391), .Z(n4421) );
  CNR2X1 U6847 ( .A(\m1.need ), .B(\m2.need ), .Z(n3392) );
  CND2X1 U6848 ( .A(n3392), .B(\m5.need ), .Z(n3393) );
  CNR2X1 U6849 ( .A(\m3.need ), .B(\m4.need ), .Z(n3398) );
  COND1XL U6850 ( .A(\m0.need ), .B(n3393), .C(n3398), .Z(n3394) );
  CNR2XL U6851 ( .A(n3394), .B(\m6.need ), .Z(n3395) );
  CNR3XL U6852 ( .A(n1846), .B(n3401), .C(n3395), .Z(n3396) );
  COND1XL U6853 ( .A(n3402), .B(n3396), .C(n5518), .Z(\nx_st[2] ) );
  CNR3XL U6854 ( .A(\m5.need ), .B(\m1.need ), .C(\m2.need ), .Z(n3397) );
  CNR2X1 U6855 ( .A(n3397), .B(\m0.need ), .Z(n3399) );
  COND1XL U6856 ( .A(\m6.need ), .B(n3399), .C(n3398), .Z(n3400) );
  COND11XL U6857 ( .A(n3402), .B(n3401), .C(n3400), .D(n1871), .Z(n3403) );
  CIVXL U6858 ( .A(n3403), .Z(n4418) );
  CIVDX3 U6859 ( .A(n3410), .Z0(\s13.addr[13] ), .Z1(n3330) );
  CIVX12 U6860 ( .A(\s13.addr[13] ), .Z(n4259) );
  CIVX2 U6861 ( .A(n3483), .Z(n4210) );
  CNR2XL U6862 ( .A(n3406), .B(n4210), .Z(\s14.SbusIn [23]) );
  CNIVX4 U6863 ( .A(n3407), .Z(n3408) );
  CIVX12 U6864 ( .A(n3408), .Z(\s12.addr[16] ) );
  CAN2XL U6865 ( .A(\s12.addr[16] ), .B(n3479), .Z(\s12.addr [62]) );
  CIVX2 U6866 ( .A(n3464), .Z(n4285) );
  CNR2XL U6867 ( .A(n2223), .B(n4285), .Z(\s8.addr [37]) );
  CAN2XL U6868 ( .A(\s8.en ), .B(n4195), .Z(\s8.addr [26]) );
  CNR2IXL U6869 ( .B(n3473), .A(n3416), .Z(\s10.SbusIn [22]) );
  CAN2XL U6870 ( .A(\s8.addr[17] ), .B(n3409), .Z(\s8.addr [7]) );
  CAN2X1 U6871 ( .A(\s8.addr[17] ), .B(n4243), .Z(\s8.SbusIn [4]) );
  CNR2XL U6872 ( .A(n2223), .B(n4253), .Z(\s8.addr [5]) );
  CAN2X1 U6873 ( .A(\s10.addr[9] ), .B(n4190), .Z(\s10.SbusIn [1]) );
  CAN2X1 U6874 ( .A(\s10.addr[9] ), .B(n4126), .Z(\s10.SbusIn [62]) );
  CIVDX3 U6875 ( .A(n3410), .Z0(\s13.addr[18] ), .Z1(n3375) );
  CIVX12 U6876 ( .A(\s13.addr[18] ), .Z(n4258) );
  CAN2X1 U6877 ( .A(\s10.addr[9] ), .B(n3467), .Z(\s10.addr [27]) );
  CAN2X1 U6878 ( .A(\s10.addr[9] ), .B(n3461), .Z(\s10.SbusIn [55]) );
  CAN2X1 U6879 ( .A(\s10.addr[9] ), .B(n4138), .Z(\s10.SbusIn [44]) );
  CIVX2 U6880 ( .A(n3469), .Z(n4228) );
  CNR2XL U6881 ( .A(n2223), .B(n4228), .Z(\s8.SbusIn [5]) );
  CAN2X1 U6882 ( .A(\s12.addr[11] ), .B(n4242), .Z(\s12.addr [56]) );
  CIVX2 U6883 ( .A(n3480), .Z(n4194) );
  CNR2XL U6884 ( .A(n3414), .B(n4194), .Z(\s12.SbusIn [49]) );
  CAN2X1 U6885 ( .A(n5445), .B(n4177), .Z(\s5.addr [39]) );
  CAN2X1 U6886 ( .A(\s12.addr[11] ), .B(n4129), .Z(\s12.SbusIn [45]) );
  CAN2X1 U6887 ( .A(\s7.en ), .B(n4125), .Z(\s7.SbusIn [61]) );
  CIVX2 U6888 ( .A(n3481), .Z(n4302) );
  CNR2XL U6889 ( .A(n2223), .B(n4302), .Z(\s8.SbusIn [12]) );
  CAN2X1 U6890 ( .A(\s12.addr[11] ), .B(n4149), .Z(\s12.SbusIn [24]) );
  CIVX2 U6891 ( .A(n3472), .Z(n4289) );
  CNR2X2 U6892 ( .A(n3418), .B(n4289), .Z(\s8.SbusIn [46]) );
  CIVX2 U6893 ( .A(n3487), .Z(n4288) );
  CNR2XL U6894 ( .A(n3416), .B(n4288), .Z(\s10.SbusIn [16]) );
  CIVX2 U6895 ( .A(n3466), .Z(n4213) );
  CNR2XL U6896 ( .A(n3417), .B(n4213), .Z(\s11.SbusIn [52]) );
  CAN2X1 U6897 ( .A(\s11.en ), .B(n4237), .Z(\s11.SbusIn [35]) );
  CAN2X1 U6898 ( .A(\s11.addr[17] ), .B(n4137), .Z(\s11.addr [48]) );
  CAN2X1 U6899 ( .A(\s11.addr[17] ), .B(n3467), .Z(\s11.addr [27]) );
  CAN2X1 U6900 ( .A(\s11.addr[17] ), .B(n4142), .Z(\s11.SbusIn [41]) );
  CAN2X1 U6901 ( .A(\s11.addr[17] ), .B(n3482), .Z(\s11.addr [60]) );
  CAN2X1 U6902 ( .A(\s11.addr[17] ), .B(n3462), .Z(\s11.addr [22]) );
  CAN2X1 U6903 ( .A(\s11.addr[17] ), .B(n4132), .Z(\s11.SbusIn [43]) );
  CAN2X1 U6904 ( .A(\s11.addr[17] ), .B(n4128), .Z(\s11.addr [21]) );
  CAN2X1 U6905 ( .A(\s11.addr[17] ), .B(n4156), .Z(\s11.SbusIn [33]) );
  CAN2X1 U6906 ( .A(n4332), .B(n4154), .Z(\s11.SbusIn [7]) );
  CAN2X1 U6907 ( .A(\s11.addr[17] ), .B(n4150), .Z(\s11.SbusIn [20]) );
  CAN2X1 U6908 ( .A(\s11.addr[17] ), .B(n4155), .Z(\s11.addr [49]) );
  CAN2X1 U6909 ( .A(n4332), .B(n4171), .Z(\s11.SbusIn [32]) );
  CAN2X1 U6910 ( .A(\s11.addr[17] ), .B(n3461), .Z(\s11.SbusIn [55]) );
  CAN2X1 U6911 ( .A(\s11.addr[17] ), .B(n4163), .Z(\s11.SbusIn [51]) );
  CAN2X1 U6912 ( .A(n4332), .B(n4149), .Z(\s11.SbusIn [24]) );
  CAN2X1 U6913 ( .A(\s11.addr[17] ), .B(n4158), .Z(\s11.SbusIn [21]) );
  CAN2X1 U6914 ( .A(\s11.addr[17] ), .B(n3470), .Z(\s11.addr [44]) );
  CAN2X1 U6915 ( .A(n4332), .B(n4135), .Z(\s11.SbusIn [39]) );
  CAN2X1 U6916 ( .A(\s11.addr[17] ), .B(n4152), .Z(\s11.SbusIn [19]) );
  CAN2X1 U6917 ( .A(n4332), .B(n4170), .Z(\s11.SbusIn [53]) );
  CAN2X1 U6918 ( .A(n4332), .B(n4123), .Z(\s11.SbusIn [13]) );
  CAN2X1 U6919 ( .A(\s11.addr[17] ), .B(n4130), .Z(\s11.SbusIn [59]) );
  CAN2X1 U6920 ( .A(n4332), .B(n4145), .Z(\s11.SbusIn [30]) );
  CAN2X1 U6921 ( .A(\s11.addr[17] ), .B(n4116), .Z(\s11.SbusIn [8]) );
  CAN2X1 U6922 ( .A(n4332), .B(n4215), .Z(\s11.SbusIn [36]) );
  CAN2X1 U6923 ( .A(\s11.addr[17] ), .B(n4192), .Z(\s11.SbusIn [2]) );
  CAN2X1 U6924 ( .A(n4332), .B(n4232), .Z(\s11.SbusIn [38]) );
  CAN2X1 U6925 ( .A(\s11.addr[17] ), .B(n4125), .Z(\s11.SbusIn [61]) );
  CAN2X1 U6926 ( .A(n4332), .B(n4121), .Z(\s11.SbusIn [48]) );
  CAN2X1 U6927 ( .A(n4332), .B(n4243), .Z(\s11.SbusIn [4]) );
  CAN2X1 U6928 ( .A(\s11.addr[17] ), .B(n3472), .Z(\s11.SbusIn [46]) );
  CAN2X1 U6929 ( .A(\s11.addr[17] ), .B(n4144), .Z(\s11.SbusIn [42]) );
  CIVX2 U6930 ( .A(n3465), .Z(n4209) );
  CNR2XL U6931 ( .A(n3417), .B(n4209), .Z(\s11.SbusIn [11]) );
  CIVX2 U6932 ( .A(n3462), .Z(n4230) );
  CNR2X2 U6933 ( .A(n3418), .B(n4230), .Z(\s8.addr [22]) );
  CIVDX4 U6934 ( .A(n3457), .Z0(n3419), .Z1(n3377) );
  CIVX16 U6935 ( .A(n3419), .Z(n4255) );
  CNR2X1 U6936 ( .A(n4255), .B(n3447), .Z(\s2.addr [8]) );
  CAN2X1 U6937 ( .A(n4405), .B(n4166), .Z(\s5.addr [52]) );
  CAN2XL U6938 ( .A(n4405), .B(n4161), .Z(\s5.SbusIn [57]) );
  CAN2XL U6939 ( .A(\s6.en ), .B(n4190), .Z(\s6.SbusIn [1]) );
  CAN2XL U6940 ( .A(\s6.en ), .B(n4200), .Z(\s6.SbusIn [3]) );
  CAN2XL U6941 ( .A(n1844), .B(n4168), .Z(\s5.SbusIn [58]) );
  CAN2XL U6942 ( .A(\s6.en ), .B(n3469), .Z(\s6.SbusIn [5]) );
  CAN2XL U6943 ( .A(\s6.en ), .B(n4329), .Z(\s6.SbusIn [6]) );
  CAN2XL U6944 ( .A(n5445), .B(n3462), .Z(\s5.addr [22]) );
  CAN2XL U6945 ( .A(\s6.en ), .B(n4154), .Z(\s6.SbusIn [7]) );
  CAN2XL U6946 ( .A(n4405), .B(n4328), .Z(\s5.addr [25]) );
  CAN2XL U6947 ( .A(\s6.en ), .B(n3481), .Z(\s6.SbusIn [12]) );
  CAN2XL U6948 ( .A(\s6.en ), .B(n4123), .Z(\s6.SbusIn [13]) );
  CAN2XL U6949 ( .A(n4405), .B(n4134), .Z(\s5.addr [29]) );
  CAN2XL U6950 ( .A(n4405), .B(n4164), .Z(\s5.addr [50]) );
  CAN2XL U6951 ( .A(\s6.en ), .B(n3483), .Z(\s6.SbusIn [23]) );
  CAN2XL U6952 ( .A(\s6.en ), .B(n4147), .Z(\s6.SbusIn [26]) );
  CAN2XL U6953 ( .A(n4405), .B(n4151), .Z(\s5.addr [61]) );
  CAN2XL U6954 ( .A(\s6.en ), .B(n4132), .Z(\s6.SbusIn [43]) );
  CAN2X1 U6955 ( .A(n3420), .B(\m3.addrM64 [63]), .Z(n3421) );
  CND2X1 U6956 ( .A(n3434), .B(\m0.addrM64 [63]), .Z(n3423) );
  CNR2IX1 U6957 ( .B(\m5.addrM64 [63]), .A(n3432), .Z(n3422) );
  CNR2IX1 U6958 ( .B(n3423), .A(n3422), .Z(n3428) );
  CAN2XL U6959 ( .A(n3424), .B(\m4.addrM64 [63]), .Z(n3425) );
  CNR2X1 U6960 ( .A(n3426), .B(n3425), .Z(n3427) );
  CND3X2 U6961 ( .A(n3429), .B(n3428), .C(n3427), .Z(n4140) );
  CAN2XL U6962 ( .A(n1844), .B(n4140), .Z(\s5.addr [63]) );
  CAN2XL U6963 ( .A(\s6.en ), .B(n4121), .Z(\s6.SbusIn [48]) );
  CAN2XL U6964 ( .A(\s6.en ), .B(n4175), .Z(\s6.SbusIn [54]) );
  CAN2XL U6965 ( .A(\s6.en ), .B(n4156), .Z(\s6.SbusIn [33]) );
  CAN2XL U6966 ( .A(\s6.en ), .B(n4143), .Z(\s6.SbusIn [40]) );
  CAN2XL U6967 ( .A(\s6.en ), .B(n4142), .Z(\s6.SbusIn [41]) );
  CAN2XL U6968 ( .A(\s6.en ), .B(n4178), .Z(\s6.SbusIn [34]) );
  CAN2XL U6969 ( .A(\s6.en ), .B(n4196), .Z(\s6.SbusIn [37]) );
  CAN2XL U6970 ( .A(\s6.en ), .B(n4232), .Z(\s6.SbusIn [38]) );
  CAN2XL U6971 ( .A(\s6.en ), .B(n4168), .Z(\s6.SbusIn [58]) );
  CAN2XL U6972 ( .A(\s6.en ), .B(n4116), .Z(\s6.SbusIn [8]) );
  CAN2XL U6973 ( .A(\s6.en ), .B(n4199), .Z(\s6.addr [24]) );
  CANR2X1 U6974 ( .A(n3431), .B(\m1.addrM64 [30]), .C(\m3.addrM64 [30]), .D(
        n3430), .Z(n3444) );
  CNR2IX1 U6975 ( .B(\m5.addrM64 [30]), .A(n3432), .Z(n3433) );
  CANR1X1 U6976 ( .A(n3434), .B(\m0.addrM64 [30]), .C(n3433), .Z(n3443) );
  CND2X1 U6977 ( .A(n3435), .B(\m6.addrM64 [30]), .Z(n3438) );
  CND2X1 U6978 ( .A(n3436), .B(\m2.addrM64 [30]), .Z(n3437) );
  CND2X1 U6979 ( .A(n3438), .B(n3437), .Z(n3441) );
  CNR2IX1 U6980 ( .B(\m4.addrM64 [30]), .A(n3439), .Z(n3440) );
  CNR2X1 U6981 ( .A(n3441), .B(n3440), .Z(n3442) );
  CND3X2 U6982 ( .A(n3444), .B(n3443), .C(n3442), .Z(n4176) );
  CAN2XL U6983 ( .A(\s6.en ), .B(n4176), .Z(\s6.addr [30]) );
  CAN2XL U6984 ( .A(\s6.en ), .B(n4180), .Z(\s6.SbusIn [18]) );
  CAN2XL U6985 ( .A(\s6.en ), .B(n4141), .Z(\s6.SbusIn [25]) );
  CAN2XL U6986 ( .A(\s6.en ), .B(n4160), .Z(\s6.addr [31]) );
  CAN2XL U6987 ( .A(\s6.en ), .B(n4145), .Z(\s6.SbusIn [30]) );
  CAN2X1 U6988 ( .A(n4405), .B(n4148), .Z(\s5.addr [54]) );
  CAN2XL U6989 ( .A(\s6.en ), .B(n4144), .Z(\s6.SbusIn [42]) );
  CNR2X1 U6990 ( .A(n3445), .B(n4254), .Z(\s4.addr [4]) );
  CAN2XL U6991 ( .A(\s6.en ), .B(n3472), .Z(\s6.SbusIn [46]) );
  CAN2XL U6992 ( .A(\s6.en ), .B(n3471), .Z(\s6.addr [41]) );
  CAN2XL U6993 ( .A(\s6.en ), .B(n4139), .Z(\s6.SbusIn [47]) );
  CAN2XL U6994 ( .A(\s6.en ), .B(n3461), .Z(\s6.SbusIn [55]) );
  CAN2XL U6995 ( .A(\s6.en ), .B(n4166), .Z(\s6.addr [52]) );
  CAN2XL U6996 ( .A(\s6.en ), .B(n4159), .Z(\s6.SbusIn [56]) );
  CAN2XL U6997 ( .A(\s6.en ), .B(n4161), .Z(\s6.SbusIn [57]) );
  CAN2XL U6998 ( .A(\s6.en ), .B(n4202), .Z(\s6.addr [58]) );
  CIVX2 U6999 ( .A(n3479), .Z(n4250) );
  CNR2X1 U7000 ( .A(n4317), .B(n4250), .Z(\s0.addr [62]) );
  CAN2XL U7001 ( .A(\s6.en ), .B(n4120), .Z(\s6.SbusIn [63]) );
  CAN2XL U7002 ( .A(\s1.addr[17] ), .B(n4180), .Z(\s1.SbusIn [18]) );
  CAN2XL U7003 ( .A(\s6.en ), .B(n4207), .Z(\s6.addr [57]) );
  CAN2XL U7004 ( .A(\s6.en ), .B(n3479), .Z(\s6.addr [62]) );
  CAN2XL U7005 ( .A(\s6.en ), .B(n4151), .Z(\s6.addr [61]) );
  CAN2XL U7006 ( .A(\s1.addr[17] ), .B(n3461), .Z(\s1.SbusIn [55]) );
  CAN2XL U7007 ( .A(\s6.en ), .B(n4140), .Z(\s6.addr [63]) );
  CAN2X1 U7008 ( .A(\s3.addr[14] ), .B(n4193), .Z(\s3.SbusIn [9]) );
  CAN2XL U7009 ( .A(\s1.addr[17] ), .B(n4155), .Z(\s1.addr [49]) );
  CAN2XL U7010 ( .A(\s1.addr[17] ), .B(n3476), .Z(\s1.addr [5]) );
  CIVX2 U7011 ( .A(n4337), .Z(n4272) );
  CNR2X1 U7012 ( .A(n3446), .B(n4272), .Z(\s1.addr [0]) );
  CAN2X1 U7013 ( .A(\s3.addr[14] ), .B(n4123), .Z(\s3.SbusIn [13]) );
  CAN2XL U7014 ( .A(\s14.addr[18] ), .B(n4329), .Z(\s14.SbusIn [6]) );
  CAN2XL U7015 ( .A(\s14.addr[17] ), .B(n4115), .Z(\s14.SbusIn [10]) );
  CAN2X1 U7016 ( .A(\s3.addr[14] ), .B(n4140), .Z(\s3.addr [63]) );
  CAN2XL U7017 ( .A(\s14.addr[18] ), .B(n3474), .Z(\s14.SbusIn [14]) );
  CAN2X1 U7018 ( .A(\s3.addr[14] ), .B(n4130), .Z(\s3.SbusIn [59]) );
  CAN2XL U7019 ( .A(\s14.addr[17] ), .B(n4193), .Z(\s14.SbusIn [9]) );
  CAN2XL U7020 ( .A(\s14.addr[18] ), .B(n4169), .Z(\s14.SbusIn [15]) );
  CAN2XL U7021 ( .A(\s14.addr[17] ), .B(n4123), .Z(\s14.SbusIn [13]) );
  CAN2XL U7022 ( .A(\s14.addr[18] ), .B(n4152), .Z(\s14.SbusIn [19]) );
  CAN2XL U7023 ( .A(\s14.addr[17] ), .B(n3481), .Z(\s14.SbusIn [12]) );
  CAN2XL U7024 ( .A(\s14.addr[18] ), .B(n4150), .Z(\s14.SbusIn [20]) );
  CAN2XL U7025 ( .A(\s14.addr [11]), .B(n4190), .Z(\s14.SbusIn [1]) );
  CAN2X1 U7026 ( .A(\s10.addr[9] ), .B(n3469), .Z(\s10.SbusIn [5]) );
  CAN2XL U7027 ( .A(\s14.addr[18] ), .B(n4158), .Z(\s14.SbusIn [21]) );
  CAN2XL U7028 ( .A(\s14.addr[17] ), .B(n4145), .Z(\s14.SbusIn [30]) );
  CNR2X1 U7029 ( .A(n4259), .B(n3447), .Z(\s13.addr [8]) );
  CNR2X1 U7030 ( .A(n4259), .B(n3448), .Z(\s13.addr [11]) );
  CNR2X1 U7031 ( .A(n4259), .B(n3468), .Z(\s13.addr [1]) );
  CAN2XL U7032 ( .A(\s14.addr[18] ), .B(n4149), .Z(\s14.SbusIn [24]) );
  CAN2XL U7033 ( .A(\s14.addr[17] ), .B(n4171), .Z(\s14.SbusIn [32]) );
  CAN2XL U7034 ( .A(\s14.addr[18] ), .B(n4141), .Z(\s14.SbusIn [25]) );
  CAN2XL U7035 ( .A(\s14.addr[17] ), .B(n4215), .Z(\s14.SbusIn [36]) );
  CAN2XL U7036 ( .A(\s14.addr [11]), .B(n3469), .Z(\s14.SbusIn [5]) );
  CAN2XL U7037 ( .A(\s14.addr [11]), .B(n4172), .Z(\s14.SbusIn [17]) );
  CAN2XL U7038 ( .A(\s14.addr[18] ), .B(n4147), .Z(\s14.SbusIn [26]) );
  CAN2XL U7039 ( .A(\s14.addr[17] ), .B(n4143), .Z(\s14.SbusIn [40]) );
  CAN2XL U7040 ( .A(\s14.addr[18] ), .B(n3460), .Z(\s14.SbusIn [27]) );
  CAN2XL U7041 ( .A(\s14.addr[17] ), .B(n4144), .Z(\s14.SbusIn [42]) );
  CAN2XL U7042 ( .A(\s14.addr[18] ), .B(n4117), .Z(\s14.SbusIn [28]) );
  CAN2XL U7043 ( .A(\s14.addr [11]), .B(n3472), .Z(\s14.SbusIn [46]) );
  CAN2XL U7044 ( .A(\s14.addr[17] ), .B(n4129), .Z(\s14.SbusIn [45]) );
  CAN2XL U7045 ( .A(\s14.addr[18] ), .B(n4197), .Z(\s14.SbusIn [29]) );
  CAN2XL U7046 ( .A(\s14.addr [11]), .B(n3465), .Z(\s14.SbusIn [11]) );
  CAN2XL U7047 ( .A(\s14.addr[17] ), .B(n4127), .Z(\s14.SbusIn [50]) );
  CAN2XL U7048 ( .A(\s9.en ), .B(n4200), .Z(\s9.SbusIn [3]) );
  CIVX2 U7049 ( .A(n3486), .Z(n4312) );
  CNR2X1 U7050 ( .A(n3451), .B(n4312), .Z(\s7.addr [40]) );
  CAN2X1 U7051 ( .A(\s10.addr [17]), .B(n4192), .Z(\s10.SbusIn [2]) );
  CAN2XL U7052 ( .A(\s14.addr[18] ), .B(n4178), .Z(\s14.SbusIn [34]) );
  CAN2X1 U7053 ( .A(\s10.addr [17]), .B(n4329), .Z(\s10.SbusIn [6]) );
  CAN2XL U7054 ( .A(\s14.addr[17] ), .B(n4139), .Z(\s14.SbusIn [47]) );
  CAN2XL U7055 ( .A(\s14.addr [11]), .B(n4243), .Z(\s14.SbusIn [4]) );
  CAN2X1 U7056 ( .A(\s10.addr [17]), .B(n3465), .Z(\s10.SbusIn [11]) );
  CAN2XL U7057 ( .A(\s14.addr[18] ), .B(n4138), .Z(\s14.SbusIn [44]) );
  CAN2X1 U7058 ( .A(\s10.addr [17]), .B(n4169), .Z(\s10.SbusIn [15]) );
  CAN2XL U7059 ( .A(n4405), .B(n4118), .Z(\s5.addr [23]) );
  CAN2XL U7060 ( .A(\s14.addr [11]), .B(n4156), .Z(\s14.SbusIn [33]) );
  CAN2X1 U7061 ( .A(\s10.addr [17]), .B(n4158), .Z(\s10.SbusIn [21]) );
  CAN2XL U7062 ( .A(\s14.addr[17] ), .B(n3466), .Z(\s14.SbusIn [52]) );
  CAN2XL U7063 ( .A(n5590), .B(n4185), .Z(\s9.SbusIn [0]) );
  CAN2X1 U7064 ( .A(\s10.addr [17]), .B(n4152), .Z(\s10.SbusIn [19]) );
  CAN2XL U7065 ( .A(\s14.addr[18] ), .B(n4121), .Z(\s14.SbusIn [48]) );
  CAN2XL U7066 ( .A(\s9.addr[7] ), .B(n4141), .Z(\s9.SbusIn [25]) );
  CAN2X1 U7067 ( .A(\s10.addr [17]), .B(n4144), .Z(\s10.SbusIn [42]) );
  CAN2XL U7068 ( .A(\s14.addr[17] ), .B(n3479), .Z(\s14.addr [62]) );
  CAN2XL U7069 ( .A(\s9.en ), .B(n4243), .Z(\s9.SbusIn [4]) );
  CAN2XL U7070 ( .A(\s9.addr[7] ), .B(n4116), .Z(\s9.SbusIn [8]) );
  CAN2XL U7071 ( .A(\s9.addr[8] ), .B(n4121), .Z(\s9.SbusIn [48]) );
  CAN2XL U7072 ( .A(\s9.addr[8] ), .B(n4115), .Z(\s9.SbusIn [10]) );
  CAN2XL U7073 ( .A(\s9.addr[16] ), .B(n3474), .Z(\s9.SbusIn [14]) );
  CAN2XL U7074 ( .A(\s9.addr[16] ), .B(n3483), .Z(\s9.SbusIn [23]) );
  CAN2XL U7075 ( .A(\s3.addr[14] ), .B(n4115), .Z(\s3.SbusIn [10]) );
  CNIVX2 U7076 ( .A(n3449), .Z(n3450) );
  CNR2X1 U7077 ( .A(n3450), .B(n4254), .Z(\s3.addr [4]) );
  CIVX2 U7078 ( .A(n3460), .Z(n4212) );
  CNR2X1 U7079 ( .A(n3450), .B(n4212), .Z(\s3.SbusIn [27]) );
  CIVX2 U7080 ( .A(n3461), .Z(n4308) );
  CNR2X1 U7081 ( .A(n3450), .B(n4308), .Z(\s3.SbusIn [55]) );
  CAN2X1 U7082 ( .A(\s10.addr [17]), .B(n3483), .Z(\s10.SbusIn [23]) );
  CAN2XL U7083 ( .A(n4405), .B(n4180), .Z(\s5.SbusIn [18]) );
  CAN2XL U7084 ( .A(\s14.addr[18] ), .B(n4125), .Z(\s14.SbusIn [61]) );
  CAN2X1 U7085 ( .A(\s10.addr [17]), .B(n4149), .Z(\s10.SbusIn [24]) );
  CAN2XL U7086 ( .A(\s14.addr [11]), .B(n4135), .Z(\s14.SbusIn [39]) );
  CAN2XL U7087 ( .A(\s9.addr[7] ), .B(n3465), .Z(\s9.SbusIn [11]) );
  CAN2X1 U7088 ( .A(\s10.addr [17]), .B(n4119), .Z(\s10.SbusIn [31]) );
  CAN2XL U7089 ( .A(\s14.addr[17] ), .B(n4175), .Z(\s14.SbusIn [54]) );
  CAN2XL U7090 ( .A(\s9.addr[7] ), .B(n4237), .Z(\s9.SbusIn [35]) );
  CAN2X1 U7091 ( .A(\s10.addr [17]), .B(n4196), .Z(\s10.SbusIn [37]) );
  CAN2XL U7092 ( .A(\s14.addr [11]), .B(n3473), .Z(\s14.SbusIn [22]) );
  CAN2XL U7093 ( .A(\s14.addr[18] ), .B(n3476), .Z(\s14.addr [5]) );
  CAN2X1 U7094 ( .A(\s10.addr [17]), .B(n4143), .Z(\s10.SbusIn [40]) );
  CAN2XL U7095 ( .A(\s9.addr[8] ), .B(n4123), .Z(\s9.SbusIn [13]) );
  CAN2XL U7096 ( .A(\s9.addr[8] ), .B(n4190), .Z(\s9.SbusIn [1]) );
  CAN2XL U7097 ( .A(\s14.addr[17] ), .B(n3461), .Z(\s14.SbusIn [55]) );
  CAN2X1 U7098 ( .A(\s10.addr [17]), .B(n4142), .Z(\s10.SbusIn [41]) );
  CAN2XL U7099 ( .A(n1844), .B(n4159), .Z(\s5.SbusIn [56]) );
  CAN2XL U7100 ( .A(\s14.addr[18] ), .B(n4331), .Z(\s14.addr [20]) );
  CAN2X1 U7101 ( .A(\s10.addr [17]), .B(n4129), .Z(\s10.SbusIn [45]) );
  CAN2XL U7102 ( .A(\s9.addr[16] ), .B(n3460), .Z(\s9.SbusIn [27]) );
  CAN2XL U7103 ( .A(\s14.addr [11]), .B(n4161), .Z(\s14.SbusIn [57]) );
  CAN2XL U7104 ( .A(\s14.addr[17] ), .B(n4159), .Z(\s14.SbusIn [56]) );
  CAN2XL U7105 ( .A(\s14.addr[18] ), .B(n4128), .Z(\s14.addr [21]) );
  CAN2XL U7106 ( .A(n5445), .B(n4174), .Z(\s5.addr [53]) );
  CAN2XL U7107 ( .A(\s9.addr[16] ), .B(n4331), .Z(\s9.addr [20]) );
  CAN2XL U7108 ( .A(\s10.addr [17]), .B(n4139), .Z(\s10.SbusIn [47]) );
  CAN2XL U7109 ( .A(\s14.addr [11]), .B(n4167), .Z(\s14.SbusIn [60]) );
  CAN2XL U7110 ( .A(\s9.addr[8] ), .B(n4144), .Z(\s9.SbusIn [42]) );
  CAN2X1 U7111 ( .A(\s10.addr [17]), .B(n3472), .Z(\s10.SbusIn [46]) );
  CAN2XL U7112 ( .A(\s14.addr[17] ), .B(n4168), .Z(\s14.SbusIn [58]) );
  CAN2XL U7113 ( .A(\s14.addr[18] ), .B(n3462), .Z(\s14.addr [22]) );
  CAN2X1 U7114 ( .A(\s10.addr [17]), .B(n3480), .Z(\s10.SbusIn [49]) );
  CAN2XL U7115 ( .A(\s9.en ), .B(n4232), .Z(\s9.SbusIn [38]) );
  CAN2X1 U7116 ( .A(\s10.addr [17]), .B(n4163), .Z(\s10.SbusIn [51]) );
  CAN2XL U7117 ( .A(\s9.addr[16] ), .B(n4135), .Z(\s9.SbusIn [39]) );
  CAN2XL U7118 ( .A(\s14.addr[17] ), .B(n4130), .Z(\s14.SbusIn [59]) );
  CAN2X1 U7119 ( .A(\s10.addr [17]), .B(n4127), .Z(\s10.SbusIn [50]) );
  CAN2XL U7120 ( .A(\s14.addr[18] ), .B(n3467), .Z(\s14.addr [27]) );
  CAN2XL U7121 ( .A(\s14.addr [11]), .B(n4199), .Z(\s14.addr [24]) );
  CAN2XL U7122 ( .A(n5590), .B(n4127), .Z(\s9.SbusIn [50]) );
  CAN2XL U7123 ( .A(\s3.addr[14] ), .B(n4120), .Z(\s3.SbusIn [63]) );
  CAN2XL U7124 ( .A(n5590), .B(n4330), .Z(\s9.addr [2]) );
  CAN2XL U7125 ( .A(\s14.addr[17] ), .B(n4120), .Z(\s14.SbusIn [63]) );
  CAN2XL U7126 ( .A(\s14.addr [11]), .B(n4196), .Z(\s14.SbusIn [37]) );
  CAN2XL U7127 ( .A(\s14.addr[18] ), .B(n4133), .Z(\s14.addr [28]) );
  CAN2XL U7128 ( .A(\s3.addr[9] ), .B(n3473), .Z(\s3.SbusIn [22]) );
  CAN2XL U7129 ( .A(\s3.addr [18]), .B(n4121), .Z(\s3.SbusIn [48]) );
  CAN2XL U7130 ( .A(\s3.addr[9] ), .B(n3467), .Z(\s3.addr [27]) );
  CAN2XL U7131 ( .A(\s10.addr [17]), .B(n4155), .Z(\s10.addr [49]) );
  CAN2X1 U7132 ( .A(\s10.addr [17]), .B(n4130), .Z(\s10.SbusIn [59]) );
  CAN2XL U7133 ( .A(\s9.en ), .B(n3480), .Z(\s9.SbusIn [49]) );
  CAN2XL U7134 ( .A(\s9.addr[8] ), .B(n4172), .Z(\s9.SbusIn [17]) );
  CAN2XL U7135 ( .A(\s14.addr[17] ), .B(n4330), .Z(\s14.addr [2]) );
  CAN2X1 U7136 ( .A(\s10.addr [17]), .B(n4120), .Z(\s10.SbusIn [63]) );
  CAN2XL U7137 ( .A(\s14.addr[18] ), .B(n4134), .Z(\s14.addr [29]) );
  CAN2XL U7138 ( .A(\s3.addr[14] ), .B(n4173), .Z(\s3.addr [35]) );
  CAN2XL U7139 ( .A(\s9.addr[7] ), .B(n4168), .Z(\s9.SbusIn [58]) );
  CAN2XL U7140 ( .A(\s14.addr[17] ), .B(n4164), .Z(\s14.addr [50]) );
  CAN2XL U7141 ( .A(\s3.addr [18]), .B(n4243), .Z(\s3.SbusIn [4]) );
  CAN2XL U7142 ( .A(\s14.addr[18] ), .B(n4176), .Z(\s14.addr [30]) );
  CAN2XL U7143 ( .A(\s14.addr[17] ), .B(n3464), .Z(\s14.addr [37]) );
  CAN2XL U7144 ( .A(\s10.addr [17]), .B(n3476), .Z(\s10.addr [5]) );
  CAN2XL U7145 ( .A(\s9.addr[16] ), .B(n3476), .Z(\s9.addr [5]) );
  CAN2XL U7146 ( .A(\s14.addr [11]), .B(n4232), .Z(\s14.SbusIn [38]) );
  CAN2XL U7147 ( .A(\s3.addr[9] ), .B(n3465), .Z(\s3.SbusIn [11]) );
  CAN2XL U7148 ( .A(\s3.addr[9] ), .B(n4126), .Z(\s3.SbusIn [62]) );
  CAN2XL U7149 ( .A(\s3.addr [18]), .B(n4330), .Z(\s3.addr [2]) );
  CAN2X1 U7150 ( .A(\s10.addr [17]), .B(n4199), .Z(\s10.addr [24]) );
  CAN2XL U7151 ( .A(\s9.addr[8] ), .B(n3466), .Z(\s9.SbusIn [52]) );
  CAN2XL U7152 ( .A(\s14.addr[18] ), .B(n4160), .Z(\s14.addr [31]) );
  CAN2X1 U7153 ( .A(\s10.addr [17]), .B(n4179), .Z(\s10.addr [33]) );
  CAN2XL U7154 ( .A(\s14.addr[17] ), .B(n4165), .Z(\s14.addr [51]) );
  CAN2XL U7155 ( .A(\s9.addr[7] ), .B(n4150), .Z(\s9.SbusIn [20]) );
  CAN2X1 U7156 ( .A(\s10.addr [17]), .B(n3471), .Z(\s10.addr [41]) );
  CAN2XL U7157 ( .A(\s3.addr[14] ), .B(n4133), .Z(\s3.addr [28]) );
  CAN2XL U7158 ( .A(\s9.addr[16] ), .B(n4159), .Z(\s9.SbusIn [56]) );
  CAN2X1 U7159 ( .A(\s10.addr [17]), .B(n4122), .Z(\s10.addr [43]) );
  CAN2XL U7160 ( .A(\s14.addr[18] ), .B(n4157), .Z(\s14.addr [32]) );
  CAN2XL U7161 ( .A(\s14.addr[17] ), .B(n4140), .Z(\s14.addr [63]) );
  CAN2X1 U7162 ( .A(\s10.addr [17]), .B(n4201), .Z(\s10.addr [55]) );
  CAN2XL U7163 ( .A(\s14.addr [11]), .B(n4155), .Z(\s14.addr [49]) );
  CAN2XL U7164 ( .A(\s3.addr [18]), .B(n3477), .Z(\s3.addr [59]) );
  CAN2XL U7165 ( .A(\s4.addr[14] ), .B(n4330), .Z(\s4.addr [2]) );
  CAN2X1 U7166 ( .A(\s10.addr [17]), .B(n4207), .Z(\s10.addr [57]) );
  CAN2XL U7167 ( .A(\s9.addr[7] ), .B(n4160), .Z(\s9.addr [31]) );
  CAN2XL U7168 ( .A(\s9.addr[8] ), .B(n4118), .Z(\s9.addr [23]) );
  CAN2XL U7169 ( .A(\s3.addr[14] ), .B(n4329), .Z(\s3.SbusIn [6]) );
  CAN2X1 U7170 ( .A(\s7.addr[19] ), .B(n4201), .Z(\s7.addr [55]) );
  CAN2X1 U7171 ( .A(\s7.en ), .B(n4176), .Z(\s7.addr [30]) );
  CAN2X1 U7172 ( .A(n4336), .B(n4333), .Z(\s7.addr [3]) );
  CAN2XL U7173 ( .A(\s14.addr [11]), .B(n4170), .Z(\s14.SbusIn [53]) );
  CAN2XL U7174 ( .A(\s3.addr[9] ), .B(n3481), .Z(\s3.SbusIn [12]) );
  CAN2XL U7175 ( .A(\s3.addr [18]), .B(n4167), .Z(\s3.SbusIn [60]) );
  CAN2XL U7176 ( .A(\s3.addr[9] ), .B(n4331), .Z(\s3.addr [20]) );
  CAN2XL U7177 ( .A(\s14.addr[18] ), .B(n4177), .Z(\s14.addr [39]) );
  CAN2XL U7178 ( .A(\s3.addr[14] ), .B(n4165), .Z(\s3.addr [51]) );
  CAN2X1 U7179 ( .A(\s7.addr[16] ), .B(n4163), .Z(\s7.SbusIn [51]) );
  CAN2XL U7180 ( .A(\s9.addr[8] ), .B(n4130), .Z(\s9.SbusIn [59]) );
  CAN2XL U7181 ( .A(\s9.addr[16] ), .B(n3473), .Z(\s9.SbusIn [22]) );
  CAN2XL U7182 ( .A(\s14.addr[18] ), .B(n3486), .Z(\s14.addr [40]) );
  CAN2X1 U7183 ( .A(n4336), .B(n3479), .Z(\s7.addr [62]) );
  CAN2XL U7184 ( .A(\s9.addr[16] ), .B(n4124), .Z(\s9.addr [36]) );
  CAN2XL U7185 ( .A(\s14.addr [11]), .B(n4118), .Z(\s14.addr [23]) );
  CAN2XL U7186 ( .A(\s3.addr [18]), .B(n4116), .Z(\s3.SbusIn [8]) );
  CAN2X1 U7187 ( .A(\s7.en ), .B(n4328), .Z(\s7.addr [25]) );
  CAN2XL U7188 ( .A(\s14.addr[18] ), .B(n3471), .Z(\s14.addr [41]) );
  CAN2XL U7189 ( .A(\s9.addr[7] ), .B(n4157), .Z(\s9.addr [32]) );
  CAN2XL U7190 ( .A(\s14.addr [11]), .B(n4195), .Z(\s14.addr [26]) );
  CAN2XL U7191 ( .A(\s3.addr [18]), .B(n4153), .Z(\s3.addr [42]) );
  CAN2XL U7192 ( .A(\s3.addr[9] ), .B(n4162), .Z(\s3.addr [45]) );
  CAN2XL U7193 ( .A(\s3.addr[9] ), .B(n4174), .Z(\s3.addr [53]) );
  CAN2XL U7194 ( .A(\s3.addr[14] ), .B(n4169), .Z(\s3.SbusIn [15]) );
  CAN2XL U7195 ( .A(\s9.addr[7] ), .B(n4126), .Z(\s9.SbusIn [62]) );
  CAN2XL U7196 ( .A(\s14.addr[18] ), .B(n4166), .Z(\s14.addr [52]) );
  CAN2XL U7197 ( .A(\s9.addr[8] ), .B(n4163), .Z(\s9.SbusIn [51]) );
  CAN2XL U7198 ( .A(n5590), .B(n4131), .Z(\s9.addr [34]) );
  CAN2XL U7199 ( .A(\s14.addr[18] ), .B(n4174), .Z(\s14.addr [53]) );
  CAN2XL U7200 ( .A(\s14.addr [11]), .B(n4328), .Z(\s14.addr [25]) );
  CAN2XL U7201 ( .A(\s3.addr [18]), .B(n4138), .Z(\s3.SbusIn [44]) );
  CAN2X1 U7202 ( .A(\s7.addr[16] ), .B(n4151), .Z(\s7.addr [61]) );
  CAN2XL U7203 ( .A(\s9.en ), .B(n4173), .Z(\s9.addr [35]) );
  CAN2XL U7204 ( .A(\s9.addr[16] ), .B(n4134), .Z(\s9.addr [29]) );
  CAN2XL U7205 ( .A(\s14.addr [11]), .B(n3456), .Z(\s14.addr [7]) );
  CAN2XL U7206 ( .A(\s3.addr[9] ), .B(n4215), .Z(\s3.SbusIn [36]) );
  CAN2XL U7207 ( .A(\s3.addr [18]), .B(n4122), .Z(\s3.addr [43]) );
  CAN2XL U7208 ( .A(\s3.addr[9] ), .B(n4146), .Z(\s3.addr [47]) );
  CAN2XL U7209 ( .A(\s14.addr[18] ), .B(n4148), .Z(\s14.addr [54]) );
  CAN2XL U7210 ( .A(\s3.addr[14] ), .B(n4175), .Z(\s3.SbusIn [54]) );
  CAN2XL U7211 ( .A(\s9.en ), .B(n4120), .Z(\s9.SbusIn [63]) );
  CAN2XL U7212 ( .A(\s9.addr[8] ), .B(n3464), .Z(\s9.addr [37]) );
  CAN2XL U7213 ( .A(\s14.addr[18] ), .B(n4207), .Z(\s14.addr [57]) );
  CAN2XL U7214 ( .A(\s14.addr [11]), .B(n4204), .Z(\s14.addr [38]) );
  CAN2XL U7215 ( .A(\s14.addr[18] ), .B(n4202), .Z(\s14.addr [58]) );
  CAN2XL U7216 ( .A(\s1.addr[17] ), .B(n3460), .Z(\s1.SbusIn [27]) );
  CAN2XL U7217 ( .A(\s3.addr[9] ), .B(n4168), .Z(\s3.SbusIn [58]) );
  CAN2XL U7218 ( .A(\s3.addr [18]), .B(n4137), .Z(\s3.addr [48]) );
  CAN2XL U7219 ( .A(\s3.addr[14] ), .B(n4156), .Z(\s3.SbusIn [33]) );
  CAN2XL U7220 ( .A(\s9.addr[16] ), .B(n3471), .Z(\s9.addr [41]) );
  CAN2XL U7221 ( .A(\s14.addr[18] ), .B(n3477), .Z(\s14.addr [59]) );
  CAN2XL U7222 ( .A(n5590), .B(n4133), .Z(\s9.addr [28]) );
  CAN2XL U7223 ( .A(\s14.addr[18] ), .B(n3482), .Z(\s14.addr [60]) );
  CAN2XL U7224 ( .A(\s9.addr[7] ), .B(n3469), .Z(\s9.SbusIn [5]) );
  CAN2XL U7225 ( .A(n5590), .B(n4329), .Z(\s9.SbusIn [6]) );
  CAN2XL U7226 ( .A(\s1.addr[17] ), .B(n4156), .Z(\s1.SbusIn [33]) );
  CAN2XL U7227 ( .A(\s3.addr [18]), .B(n4148), .Z(\s3.addr [54]) );
  CAN2XL U7228 ( .A(\s9.addr[7] ), .B(n4179), .Z(\s9.addr [33]) );
  CAN2XL U7229 ( .A(\s9.en ), .B(n4193), .Z(\s9.SbusIn [9]) );
  CAN2XL U7230 ( .A(\s9.addr[8] ), .B(n4180), .Z(\s9.SbusIn [18]) );
  CAN2XL U7231 ( .A(\s1.addr[17] ), .B(n4125), .Z(\s1.SbusIn [61]) );
  CIVDX1 U7232 ( .A(n3474), .Z0(n4225) );
  CNR2X1 U7233 ( .A(n3451), .B(n4225), .Z(\s7.SbusIn [14]) );
  CAN2X1 U7234 ( .A(\s1.addr[15] ), .B(n4237), .Z(\s1.SbusIn [35]) );
  CAN2XL U7235 ( .A(\s1.addr[17] ), .B(n4330), .Z(\s1.addr [2]) );
  CAN2XL U7236 ( .A(\s12.addr[10] ), .B(n4207), .Z(\s12.addr [57]) );
  CAN2XL U7237 ( .A(\s7.addr[19] ), .B(n3465), .Z(\s7.SbusIn [11]) );
  CAN2XL U7238 ( .A(\s1.addr[15] ), .B(n4164), .Z(\s1.addr [50]) );
  CAN2XL U7239 ( .A(\s9.addr[16] ), .B(n4158), .Z(\s9.SbusIn [21]) );
  CAN2XL U7240 ( .A(\s9.addr[7] ), .B(n4145), .Z(\s9.SbusIn [30]) );
  CAN2XL U7241 ( .A(\s7.en ), .B(n4169), .Z(\s7.SbusIn [15]) );
  CAN2XL U7242 ( .A(n4336), .B(n4158), .Z(\s7.SbusIn [21]) );
  CAN2XL U7243 ( .A(\s9.addr[16] ), .B(n3481), .Z(\s9.SbusIn [12]) );
  CAN2XL U7244 ( .A(\s7.addr[16] ), .B(n3483), .Z(\s7.SbusIn [23]) );
  CAN2XL U7245 ( .A(\s9.addr[8] ), .B(n4149), .Z(\s9.SbusIn [24]) );
  CAN2XL U7246 ( .A(\s9.addr[16] ), .B(n4156), .Z(\s9.SbusIn [33]) );
  CNR2X1 U7247 ( .A(n3453), .B(n4254), .Z(\s1.addr [4]) );
  CAN2XL U7248 ( .A(\s7.addr[19] ), .B(n4149), .Z(\s7.SbusIn [24]) );
  CAN2XL U7249 ( .A(n5590), .B(n4197), .Z(\s9.SbusIn [29]) );
  CNR2X1 U7250 ( .A(n4258), .B(n4254), .Z(\s13.addr [4]) );
  CAN2XL U7251 ( .A(\s7.en ), .B(n4119), .Z(\s7.SbusIn [31]) );
  CAN2XL U7252 ( .A(\s9.addr[7] ), .B(n4215), .Z(\s9.SbusIn [36]) );
  CAN2XL U7253 ( .A(\s9.addr[8] ), .B(n4196), .Z(\s9.SbusIn [37]) );
  CAN2XL U7254 ( .A(\s7.en ), .B(n4171), .Z(\s7.SbusIn [32]) );
  CAN2XL U7255 ( .A(\s9.en ), .B(n4138), .Z(\s9.SbusIn [44]) );
  CAN2XL U7256 ( .A(\s10.en ), .B(n3466), .Z(\s10.SbusIn [52]) );
  CAN2XL U7257 ( .A(n4336), .B(n4143), .Z(\s7.SbusIn [40]) );
  CAN2XL U7258 ( .A(\s9.addr[16] ), .B(n4170), .Z(\s9.SbusIn [53]) );
  CAN2XL U7259 ( .A(\s9.en ), .B(n4177), .Z(\s9.addr [39]) );
  CAN2XL U7260 ( .A(\s7.addr[19] ), .B(n4161), .Z(\s7.SbusIn [57]) );
  CNR2X1 U7261 ( .A(n4258), .B(n3454), .Z(\s13.addr [9]) );
  CNR2X1 U7262 ( .A(n4258), .B(n3459), .Z(\s13.addr [3]) );
  CAN2XL U7263 ( .A(\s9.addr[8] ), .B(n4142), .Z(\s9.SbusIn [41]) );
  CAN2XL U7264 ( .A(\s7.addr[16] ), .B(n3480), .Z(\s7.SbusIn [49]) );
  CAN2XL U7265 ( .A(\s10.addr[9] ), .B(n4156), .Z(\s10.SbusIn [33]) );
  CAN2XL U7266 ( .A(\s1.addr[15] ), .B(n3469), .Z(\s1.SbusIn [5]) );
  CAN2XL U7267 ( .A(\s1.en ), .B(n4192), .Z(\s1.SbusIn [2]) );
  CAN2XL U7268 ( .A(\s1.addr [19]), .B(n3465), .Z(\s1.SbusIn [11]) );
  CAN2XL U7269 ( .A(n5590), .B(n4176), .Z(\s9.addr [30]) );
  CAN2XL U7270 ( .A(\s9.addr[7] ), .B(n4136), .Z(\s9.addr [46]) );
  CAN2XL U7271 ( .A(\s7.en ), .B(n4168), .Z(\s7.SbusIn [58]) );
  CAN2XL U7272 ( .A(\s9.addr[16] ), .B(n4139), .Z(\s9.SbusIn [47]) );
  CAN2XL U7273 ( .A(\s1.en ), .B(n4243), .Z(\s1.SbusIn [4]) );
  CAN2XL U7274 ( .A(\s1.addr [19]), .B(n4136), .Z(\s1.addr [46]) );
  CAN2XL U7275 ( .A(n4336), .B(n4127), .Z(\s7.SbusIn [50]) );
  CAN2XL U7276 ( .A(\s9.addr[8] ), .B(n4175), .Z(\s9.SbusIn [54]) );
  CAN2XL U7277 ( .A(\s9.addr[16] ), .B(n4204), .Z(\s9.addr [38]) );
  CAN2XL U7278 ( .A(\s1.addr [19]), .B(n3474), .Z(\s1.SbusIn [14]) );
  CAN2XL U7279 ( .A(\s1.en ), .B(n4158), .Z(\s1.SbusIn [21]) );
  CAN2XL U7280 ( .A(\s1.en ), .B(n4329), .Z(\s1.SbusIn [6]) );
  CAN2X1 U7281 ( .A(\s7.addr[16] ), .B(n4185), .Z(\s7.SbusIn [0]) );
  CAN2X1 U7282 ( .A(n4336), .B(n4192), .Z(\s7.SbusIn [2]) );
  CAN2XL U7283 ( .A(\s9.addr[7] ), .B(n4125), .Z(\s9.SbusIn [61]) );
  CAN2X1 U7284 ( .A(\s7.en ), .B(n4329), .Z(\s7.SbusIn [6]) );
  CAN2X1 U7285 ( .A(\s7.addr[19] ), .B(n3469), .Z(\s7.SbusIn [5]) );
  CAN2XL U7286 ( .A(\s1.addr [19]), .B(n4172), .Z(\s1.SbusIn [17]) );
  CAN2XL U7287 ( .A(\s1.en ), .B(n3483), .Z(\s1.SbusIn [23]) );
  CAN2XL U7288 ( .A(\s1.addr[15] ), .B(n4116), .Z(\s1.SbusIn [8]) );
  CAN2XL U7289 ( .A(\s9.addr[8] ), .B(n4153), .Z(\s9.addr [42]) );
  CAN2XL U7290 ( .A(\s9.addr[16] ), .B(n4165), .Z(\s9.addr [51]) );
  CAN2X1 U7291 ( .A(\s7.addr[16] ), .B(n4116), .Z(\s7.SbusIn [8]) );
  CAN2X1 U7292 ( .A(n4336), .B(n4147), .Z(\s7.SbusIn [26]) );
  CAN2X1 U7293 ( .A(\s7.en ), .B(n4117), .Z(\s7.SbusIn [28]) );
  CAN2XL U7294 ( .A(\s9.addr[8] ), .B(n3461), .Z(\s9.SbusIn [55]) );
  CAN2XL U7295 ( .A(\s1.addr [19]), .B(n4178), .Z(\s1.SbusIn [34]) );
  CAN2XL U7296 ( .A(\s1.en ), .B(n4232), .Z(\s1.SbusIn [38]) );
  CAN2XL U7297 ( .A(\s1.en ), .B(n4115), .Z(\s1.SbusIn [10]) );
  CAN2X1 U7298 ( .A(\s7.en ), .B(n4144), .Z(\s7.SbusIn [42]) );
  CAN2X1 U7299 ( .A(\s7.addr[19] ), .B(n4138), .Z(\s7.SbusIn [44]) );
  CAN2XL U7300 ( .A(\s9.addr[7] ), .B(n4162), .Z(\s9.addr [45]) );
  CAN2XL U7301 ( .A(n5590), .B(n4148), .Z(\s9.addr [54]) );
  CAN2XL U7302 ( .A(\s1.addr [19]), .B(n4190), .Z(\s1.SbusIn [1]) );
  CAN2XL U7303 ( .A(\s1.en ), .B(n4152), .Z(\s1.SbusIn [19]) );
  CAN2XL U7304 ( .A(\s1.addr[15] ), .B(n4185), .Z(\s1.SbusIn [0]) );
  CAN2XL U7305 ( .A(\s7.addr[16] ), .B(n4159), .Z(\s7.SbusIn [56]) );
  CAN2XL U7306 ( .A(\s7.addr[19] ), .B(n4139), .Z(\s7.SbusIn [47]) );
  CAN2X1 U7307 ( .A(\s7.en ), .B(n3466), .Z(\s7.SbusIn [52]) );
  CAN2XL U7308 ( .A(\s1.addr [19]), .B(n4196), .Z(\s1.SbusIn [37]) );
  CAN2XL U7309 ( .A(\s1.en ), .B(n4142), .Z(\s1.SbusIn [41]) );
  CAN2XL U7310 ( .A(\s1.en ), .B(n4147), .Z(\s1.SbusIn [26]) );
  CAN2XL U7311 ( .A(\s9.en ), .B(n4122), .Z(\s9.addr [43]) );
  CAN2XL U7312 ( .A(\s9.addr[8] ), .B(n4174), .Z(\s9.addr [53]) );
  CAN2X1 U7313 ( .A(\s7.addr[16] ), .B(n4167), .Z(\s7.SbusIn [60]) );
  CAN2X1 U7314 ( .A(\s7.addr[19] ), .B(n4126), .Z(\s7.SbusIn [62]) );
  CAN2XL U7315 ( .A(\s3.addr [18]), .B(n3464), .Z(\s3.addr [37]) );
  CAN2X1 U7316 ( .A(n4336), .B(n3455), .Z(\s7.addr [9]) );
  CAN2XL U7317 ( .A(\s1.addr [19]), .B(n4135), .Z(\s1.SbusIn [39]) );
  CAN2XL U7318 ( .A(\s1.en ), .B(n4132), .Z(\s1.SbusIn [43]) );
  CAN2XL U7319 ( .A(\s1.addr[15] ), .B(n4144), .Z(\s1.SbusIn [42]) );
  CAN2XL U7320 ( .A(\s12.addr[11] ), .B(n3474), .Z(\s12.SbusIn [14]) );
  CAN2XL U7321 ( .A(\s6.addr [17]), .B(n3477), .Z(\s6.addr [59]) );
  CAN2XL U7322 ( .A(\s1.addr [19]), .B(n3466), .Z(\s1.SbusIn [52]) );
  CAN2XL U7323 ( .A(\s1.en ), .B(n4130), .Z(\s1.SbusIn [59]) );
  CAN2XL U7324 ( .A(\s1.en ), .B(n4139), .Z(\s1.SbusIn [47]) );
  CAN2XL U7325 ( .A(\s1.en ), .B(n4161), .Z(\s1.SbusIn [57]) );
  CAN2XL U7326 ( .A(\s1.addr[15] ), .B(n4121), .Z(\s1.SbusIn [48]) );
  CAN2XL U7327 ( .A(\s1.en ), .B(n4168), .Z(\s1.SbusIn [58]) );
  CAN2XL U7328 ( .A(\s1.addr [19]), .B(n4133), .Z(\s1.addr [28]) );
  CAN2XL U7329 ( .A(\s1.en ), .B(n4170), .Z(\s1.SbusIn [53]) );
  CAN2XL U7330 ( .A(\s1.en ), .B(n4141), .Z(\s1.SbusIn [25]) );
  CAN2XL U7331 ( .A(\s1.addr [19]), .B(n4159), .Z(\s1.SbusIn [56]) );
  CAN2XL U7332 ( .A(\s1.addr[15] ), .B(n4169), .Z(\s1.SbusIn [15]) );
  CAN2X1 U7333 ( .A(\s12.addr[10] ), .B(n4197), .Z(\s12.SbusIn [29]) );
  CAN2X1 U7334 ( .A(\s12.addr[11] ), .B(n4117), .Z(\s12.SbusIn [28]) );
  CAN2XL U7335 ( .A(\s1.addr [19]), .B(n4134), .Z(\s1.addr [29]) );
  CAN2XL U7336 ( .A(\s1.en ), .B(n4176), .Z(\s1.addr [30]) );
  CAN2XL U7337 ( .A(\s1.en ), .B(n4120), .Z(\s1.SbusIn [63]) );
  CAN2XL U7338 ( .A(n4332), .B(n4338), .Z(\s11.addr [4]) );
  CAN2X1 U7339 ( .A(\s12.addr[10] ), .B(n4178), .Z(\s12.SbusIn [34]) );
  CAN2X1 U7340 ( .A(\s12.addr[16] ), .B(n4142), .Z(\s12.SbusIn [41]) );
  CAN2XL U7341 ( .A(\s8.addr[17] ), .B(n3460), .Z(\s8.SbusIn [27]) );
  CAN2XL U7342 ( .A(\s1.en ), .B(n3456), .Z(\s1.addr [7]) );
  CAN2XL U7343 ( .A(\s1.addr [19]), .B(n4160), .Z(\s1.addr [31]) );
  CAN2XL U7344 ( .A(\s1.addr[15] ), .B(n4118), .Z(\s1.addr [23]) );
  CAN2X1 U7345 ( .A(\s12.addr[10] ), .B(n3472), .Z(\s12.SbusIn [46]) );
  CAN2X1 U7346 ( .A(\s8.addr[15] ), .B(n4143), .Z(\s8.SbusIn [40]) );
  CAN2XL U7347 ( .A(\s1.en ), .B(n4137), .Z(\s1.addr [48]) );
  CAN2XL U7348 ( .A(\s1.addr [19]), .B(n4207), .Z(\s1.addr [57]) );
  CAN2XL U7349 ( .A(\s1.en ), .B(n3486), .Z(\s1.addr [40]) );
  CAN2XL U7350 ( .A(\s12.addr[11] ), .B(n4159), .Z(\s12.SbusIn [56]) );
  CAN2X1 U7351 ( .A(\s8.addr[15] ), .B(n4331), .Z(\s8.addr [20]) );
  CAN2XL U7352 ( .A(\s8.addr[17] ), .B(n4180), .Z(\s8.SbusIn [18]) );
  CAN2X1 U7353 ( .A(\s12.addr[11] ), .B(n4130), .Z(\s12.SbusIn [59]) );
  CAN2XL U7354 ( .A(\s8.en ), .B(n4200), .Z(\s8.SbusIn [3]) );
  CAN2X1 U7355 ( .A(\s8.addr[15] ), .B(n4149), .Z(\s8.SbusIn [24]) );
  CAN2X1 U7356 ( .A(\s12.addr[10] ), .B(n4120), .Z(\s12.SbusIn [63]) );
  CAN2XL U7357 ( .A(\s11.en ), .B(n4115), .Z(\s11.SbusIn [10]) );
  CAN2XL U7358 ( .A(\s12.addr[16] ), .B(n4118), .Z(\s12.addr [23]) );
  CAN2XL U7359 ( .A(\s8.addr[17] ), .B(n4123), .Z(\s8.SbusIn [13]) );
  CAN2X1 U7360 ( .A(\s12.addr[16] ), .B(n3464), .Z(\s12.addr [37]) );
  CAN2X1 U7361 ( .A(\s12.addr[11] ), .B(n4126), .Z(\s12.SbusIn [62]) );
  CAN2XL U7362 ( .A(\s11.en ), .B(n3474), .Z(\s11.SbusIn [14]) );
  CAN2XL U7363 ( .A(\s11.en ), .B(n4161), .Z(\s11.SbusIn [57]) );
  CAN2XL U7364 ( .A(\s12.addr[16] ), .B(n4177), .Z(\s12.addr [39]) );
  CAN2X1 U7365 ( .A(\s12.addr[10] ), .B(n4136), .Z(\s12.addr [46]) );
  CAN2X1 U7366 ( .A(\s7.addr[16] ), .B(n4154), .Z(\s7.SbusIn [7]) );
  CAN2X1 U7367 ( .A(\s12.addr[11] ), .B(n4166), .Z(\s12.addr [52]) );
  CAN2X1 U7368 ( .A(\s12.addr[16] ), .B(n4140), .Z(\s12.addr [63]) );
  CAN2XL U7369 ( .A(\s12.addr[16] ), .B(n4116), .Z(\s12.SbusIn [8]) );
  CAN2XL U7370 ( .A(n4336), .B(n3460), .Z(\s7.SbusIn [27]) );
  CAN2X1 U7371 ( .A(n4336), .B(n4130), .Z(\s7.SbusIn [59]) );
  CAN2X1 U7372 ( .A(\s7.en ), .B(n4132), .Z(\s7.SbusIn [43]) );
  CAN2XL U7373 ( .A(\s12.addr[16] ), .B(n4192), .Z(\s12.SbusIn [2]) );
  CAN2X1 U7374 ( .A(\s7.addr[19] ), .B(n4120), .Z(\s7.SbusIn [63]) );
  CAN2X1 U7375 ( .A(n4405), .B(n4202), .Z(\s5.addr [58]) );
  CAN2XL U7376 ( .A(\s12.addr[16] ), .B(n4190), .Z(\s12.SbusIn [1]) );
  CAN2XL U7377 ( .A(\s12.addr[16] ), .B(n4185), .Z(\s12.SbusIn [0]) );
  CAN2XL U7378 ( .A(\s7.en ), .B(n3476), .Z(\s7.addr [5]) );
  CAN2XL U7379 ( .A(\s11.en ), .B(n4168), .Z(\s11.SbusIn [58]) );
  CAN2XL U7380 ( .A(n4332), .B(n4120), .Z(\s11.SbusIn [63]) );
  CAN2X1 U7381 ( .A(\s7.addr[16] ), .B(n4173), .Z(\s7.addr [35]) );
  CAN2X1 U7382 ( .A(n4336), .B(n4153), .Z(\s7.addr [42]) );
  CAN2XL U7383 ( .A(\s12.addr[16] ), .B(n4243), .Z(\s12.SbusIn [4]) );
  CAN2XL U7384 ( .A(\s12.addr[16] ), .B(n4193), .Z(\s12.SbusIn [9]) );
  CAN2XL U7385 ( .A(n4332), .B(n3481), .Z(\s11.SbusIn [12]) );
  CAN2XL U7386 ( .A(\s12.addr[16] ), .B(n4154), .Z(\s12.SbusIn [7]) );
  CAN2XL U7387 ( .A(\s12.addr[16] ), .B(n3460), .Z(\s12.SbusIn [27]) );
  CAN2XL U7388 ( .A(n4332), .B(n4167), .Z(\s11.SbusIn [60]) );
  CAN2XL U7389 ( .A(\s12.addr[10] ), .B(n4172), .Z(\s12.SbusIn [17]) );
  CAN2XL U7390 ( .A(\s12.addr[16] ), .B(n4123), .Z(\s12.SbusIn [13]) );
  CAN2XL U7391 ( .A(\s12.addr[16] ), .B(n4145), .Z(\s12.SbusIn [30]) );
  CAN2XL U7392 ( .A(\s8.addr[17] ), .B(n4118), .Z(\s8.addr [23]) );
  CAN2XL U7393 ( .A(\s8.addr[17] ), .B(n3480), .Z(\s8.SbusIn [49]) );
  CAN2XL U7394 ( .A(\s8.addr[15] ), .B(n4115), .Z(\s8.SbusIn [10]) );
  CAN2XL U7395 ( .A(\s12.addr[10] ), .B(n4171), .Z(\s12.SbusIn [32]) );
  CAN2XL U7396 ( .A(\s12.addr[11] ), .B(n4141), .Z(\s12.SbusIn [25]) );
  CAN2X1 U7397 ( .A(\s12.addr[11] ), .B(n3481), .Z(\s12.SbusIn [12]) );
  CAN2XL U7398 ( .A(\s12.addr[16] ), .B(n4119), .Z(\s12.SbusIn [31]) );
  CAN2X1 U7399 ( .A(\s12.addr[11] ), .B(n4169), .Z(\s12.SbusIn [15]) );
  CAN2X1 U7400 ( .A(\s12.addr[11] ), .B(n3487), .Z(\s12.SbusIn [16]) );
  CAN2XL U7401 ( .A(\s12.addr[10] ), .B(n4127), .Z(\s12.SbusIn [50]) );
  CAN2XL U7402 ( .A(\s12.addr[16] ), .B(n4170), .Z(\s12.SbusIn [53]) );
  CAN2X1 U7403 ( .A(\s12.addr[11] ), .B(n4147), .Z(\s12.SbusIn [26]) );
  CAN2XL U7404 ( .A(\s12.addr[16] ), .B(n4125), .Z(\s12.SbusIn [61]) );
  CAN2X1 U7405 ( .A(\s12.addr[11] ), .B(n4132), .Z(\s12.SbusIn [43]) );
  CAN2XL U7406 ( .A(\s12.addr[16] ), .B(n4138), .Z(\s12.SbusIn [44]) );
  CAN2XL U7407 ( .A(\s12.addr[10] ), .B(n4215), .Z(\s12.SbusIn [36]) );
  CAN2XL U7408 ( .A(\s12.addr[16] ), .B(n4232), .Z(\s12.SbusIn [38]) );
  CAN2X1 U7409 ( .A(\s12.addr[10] ), .B(n4237), .Z(\s12.SbusIn [35]) );
  CAN2XL U7410 ( .A(\s12.addr[11] ), .B(n4156), .Z(\s12.SbusIn [33]) );
  CAN2X1 U7411 ( .A(\s12.addr[11] ), .B(n4128), .Z(\s12.addr [21]) );
  CAN2X1 U7412 ( .A(\s12.addr[11] ), .B(n3473), .Z(\s12.SbusIn [22]) );
  CAN2XL U7413 ( .A(\s10.en ), .B(n3474), .Z(\s10.SbusIn [14]) );
  CAN2XL U7414 ( .A(\s12.addr[16] ), .B(n3467), .Z(\s12.addr [27]) );
  CAN2XL U7415 ( .A(\s8.addr[17] ), .B(n4142), .Z(\s8.SbusIn [41]) );
  CAN2XL U7416 ( .A(\s12.addr[10] ), .B(n3466), .Z(\s12.SbusIn [52]) );
  CAN2X1 U7417 ( .A(\s12.addr[11] ), .B(n3462), .Z(\s12.addr [22]) );
  CAN2XL U7418 ( .A(\s12.addr[16] ), .B(n4199), .Z(\s12.addr [24]) );
  CAN2X1 U7419 ( .A(\s12.addr[11] ), .B(n4157), .Z(\s12.addr [32]) );
  CAN2X1 U7420 ( .A(\s12.addr[11] ), .B(n4173), .Z(\s12.addr [35]) );
  CAN2XL U7421 ( .A(\s11.addr[19] ), .B(n4173), .Z(\s11.addr [35]) );
  CAN2XL U7422 ( .A(\s11.addr[17] ), .B(n4124), .Z(\s11.addr [36]) );
  CAN2XL U7423 ( .A(\s11.addr[19] ), .B(n4136), .Z(\s11.addr [46]) );
  CAN2X1 U7424 ( .A(\s12.addr[11] ), .B(n4143), .Z(\s12.SbusIn [40]) );
  CAN2XL U7425 ( .A(\s12.addr[16] ), .B(n4152), .Z(\s12.SbusIn [19]) );
  CAN2XL U7426 ( .A(\s12.addr[16] ), .B(n4160), .Z(\s12.addr [31]) );
  CAN2XL U7427 ( .A(\s12.addr[10] ), .B(n4158), .Z(\s12.SbusIn [21]) );
  CAN2XL U7428 ( .A(\s12.addr[10] ), .B(n3483), .Z(\s12.SbusIn [23]) );
  CAN2XL U7429 ( .A(\s12.addr[11] ), .B(n4135), .Z(\s12.SbusIn [39]) );
  CAN2XL U7430 ( .A(\s10.en ), .B(n4180), .Z(\s10.SbusIn [18]) );
  CAN2XL U7431 ( .A(\s8.addr[17] ), .B(n4156), .Z(\s8.SbusIn [33]) );
  CAN2XL U7432 ( .A(\s12.addr[16] ), .B(n4167), .Z(\s12.SbusIn [60]) );
  CAN2XL U7433 ( .A(\s12.addr[11] ), .B(n4179), .Z(\s12.addr [33]) );
  CAN2XL U7434 ( .A(\s8.addr[17] ), .B(n4145), .Z(\s8.SbusIn [30]) );
  CAN2XL U7435 ( .A(\s12.addr[16] ), .B(n4195), .Z(\s12.addr [26]) );
  CAN2XL U7436 ( .A(\s8.addr[17] ), .B(n3483), .Z(\s8.SbusIn [23]) );
  CAN2X1 U7437 ( .A(\s10.en ), .B(n4232), .Z(\s10.SbusIn [38]) );
  CAN2XL U7438 ( .A(\s12.addr[10] ), .B(n4139), .Z(\s12.SbusIn [47]) );
  CAN2XL U7439 ( .A(\s12.addr[10] ), .B(n4150), .Z(\s12.SbusIn [20]) );
  CAN2XL U7440 ( .A(\s12.addr[11] ), .B(n4196), .Z(\s12.SbusIn [37]) );
  CAN2XL U7441 ( .A(\s7.en ), .B(n4115), .Z(\s7.SbusIn [10]) );
  CAN2X1 U7442 ( .A(\s8.addr[17] ), .B(n4172), .Z(\s8.SbusIn [17]) );
  CAN2X1 U7443 ( .A(\s8.addr[15] ), .B(n4152), .Z(\s8.SbusIn [19]) );
  CAN2X1 U7444 ( .A(\s10.en ), .B(n3456), .Z(\s10.addr [7]) );
  CAN2XL U7445 ( .A(\s8.addr[17] ), .B(n4139), .Z(\s8.SbusIn [47]) );
  CAN2XL U7446 ( .A(\s12.addr[16] ), .B(n4133), .Z(\s12.addr [28]) );
  CAN2XL U7447 ( .A(\s12.addr[16] ), .B(n4131), .Z(\s12.addr [34]) );
  CAN2XL U7448 ( .A(\s12.addr[10] ), .B(n4162), .Z(\s12.addr [45]) );
  CAN2X1 U7449 ( .A(\s10.en ), .B(n4133), .Z(\s10.addr [28]) );
  CAN2XL U7450 ( .A(\s12.addr[10] ), .B(n3461), .Z(\s12.SbusIn [55]) );
  CAN2XL U7451 ( .A(\s10.en ), .B(n4134), .Z(\s10.addr [29]) );
  CAN2XL U7452 ( .A(\s12.addr[10] ), .B(n4168), .Z(\s12.SbusIn [58]) );
  CAN2XL U7453 ( .A(\s12.addr[11] ), .B(n3471), .Z(\s12.addr [41]) );
  CAN2X1 U7454 ( .A(\s10.en ), .B(n4153), .Z(\s10.addr [42]) );
  CAN2XL U7455 ( .A(\s12.addr[16] ), .B(n4176), .Z(\s12.addr [30]) );
  CAN2XL U7456 ( .A(\s12.addr[16] ), .B(n4204), .Z(\s12.addr [38]) );
  CAN2XL U7457 ( .A(\s12.addr[11] ), .B(n4146), .Z(\s12.addr [47]) );
  CAN2X1 U7458 ( .A(\s7.en ), .B(n3473), .Z(\s7.SbusIn [22]) );
  CAN2X1 U7459 ( .A(\s10.en ), .B(n3470), .Z(\s10.addr [44]) );
  CAN2XL U7460 ( .A(\s12.addr[10] ), .B(n4161), .Z(\s12.SbusIn [57]) );
  CAN2XL U7461 ( .A(\s12.addr[10] ), .B(n4134), .Z(\s12.addr [29]) );
  CAN2XL U7462 ( .A(\s12.addr[11] ), .B(n4137), .Z(\s12.addr [48]) );
  CAN2XL U7463 ( .A(n4336), .B(n4129), .Z(\s7.SbusIn [45]) );
  CAN2X1 U7464 ( .A(\s7.en ), .B(n4197), .Z(\s7.SbusIn [29]) );
  CAN2XL U7465 ( .A(\s12.addr[16] ), .B(n4153), .Z(\s12.addr [42]) );
  CAN2XL U7466 ( .A(\s12.addr[16] ), .B(n4122), .Z(\s12.addr [43]) );
  CAN2X1 U7467 ( .A(\s10.en ), .B(n4166), .Z(\s10.addr [52]) );
  CAN2XL U7468 ( .A(\s12.addr[11] ), .B(n3477), .Z(\s12.addr [59]) );
  CAN2X1 U7469 ( .A(\s10.en ), .B(n3479), .Z(\s10.addr [62]) );
  CAN2XL U7470 ( .A(\s12.addr[10] ), .B(n4328), .Z(\s12.addr [25]) );
  CAN2XL U7471 ( .A(\s12.addr[16] ), .B(n4155), .Z(\s12.addr [49]) );
  CAN2XL U7472 ( .A(\s12.addr[10] ), .B(n4124), .Z(\s12.addr [36]) );
  CAN2XL U7473 ( .A(\s12.addr[11] ), .B(n4174), .Z(\s12.addr [53]) );
  CAN2XL U7474 ( .A(\s12.addr[16] ), .B(n4164), .Z(\s12.addr [50]) );
  CAN2XL U7475 ( .A(\s12.addr[10] ), .B(n3486), .Z(\s12.addr [40]) );
  CAN2X1 U7476 ( .A(\s10.addr [17]), .B(n3485), .Z(\s10.addr [6]) );
  CAN2XL U7477 ( .A(\s12.addr[11] ), .B(n3482), .Z(\s12.addr [60]) );
  CAN2XL U7478 ( .A(\s12.addr[16] ), .B(n4165), .Z(\s12.addr [51]) );
  CAN2XL U7479 ( .A(\s12.addr[10] ), .B(n3470), .Z(\s12.addr [44]) );
  CAN2XL U7480 ( .A(\s12.addr[10] ), .B(n4148), .Z(\s12.addr [54]) );
  CAN2XL U7481 ( .A(\s12.addr[16] ), .B(n4202), .Z(\s12.addr [58]) );
  CAN2XL U7482 ( .A(\s10.en ), .B(n4121), .Z(\s10.SbusIn [48]) );
  CAN2XL U7483 ( .A(\s12.addr[16] ), .B(n4151), .Z(\s12.addr [61]) );
  CAN2XL U7484 ( .A(\s10.addr[9] ), .B(n3460), .Z(\s10.SbusIn [27]) );
  CAN2XL U7485 ( .A(\s12.addr[10] ), .B(n3476), .Z(\s12.addr [5]) );
  CAN2XL U7486 ( .A(\s6.en ), .B(n3476), .Z(\s6.addr [5]) );
  CAN2XL U7487 ( .A(\s8.en ), .B(n4132), .Z(\s8.SbusIn [43]) );
  CAN2X1 U7488 ( .A(\s8.addr[17] ), .B(n4135), .Z(\s8.SbusIn [39]) );
  CAN2X1 U7489 ( .A(\s8.addr[15] ), .B(n4150), .Z(\s8.SbusIn [20]) );
  CAN2X1 U7490 ( .A(\s10.addr[9] ), .B(n4132), .Z(\s10.SbusIn [43]) );
  CAN2XL U7491 ( .A(\s8.addr[17] ), .B(n4144), .Z(\s8.SbusIn [42]) );
  CAN2X1 U7492 ( .A(\s8.addr[15] ), .B(n4215), .Z(\s8.SbusIn [36]) );
  CAN2X1 U7493 ( .A(\s10.addr[9] ), .B(n4237), .Z(\s10.SbusIn [35]) );
  CAN2X1 U7494 ( .A(\s10.addr[9] ), .B(n4159), .Z(\s10.SbusIn [56]) );
  CAN2X1 U7495 ( .A(\s8.addr[17] ), .B(n3466), .Z(\s8.SbusIn [52]) );
  CAN2X1 U7496 ( .A(\s8.addr[15] ), .B(n4147), .Z(\s8.SbusIn [26]) );
  CAN2X1 U7497 ( .A(\s10.addr[9] ), .B(n4160), .Z(\s10.addr [31]) );
  CAN2X1 U7498 ( .A(\s8.addr[15] ), .B(n4138), .Z(\s8.SbusIn [44]) );
  CAN2X1 U7499 ( .A(\s10.addr[9] ), .B(n4215), .Z(\s10.SbusIn [36]) );
  CAN2X1 U7500 ( .A(\s8.addr[15] ), .B(n4130), .Z(\s8.SbusIn [59]) );
  CAN2X1 U7501 ( .A(\s10.addr[9] ), .B(n4157), .Z(\s10.addr [32]) );
  CAN2XL U7502 ( .A(\s8.addr[17] ), .B(n4128), .Z(\s8.addr [21]) );
  CAN2X1 U7503 ( .A(\s8.addr[15] ), .B(n4232), .Z(\s8.SbusIn [38]) );
  CAN2X1 U7504 ( .A(\s10.addr[9] ), .B(n4170), .Z(\s10.SbusIn [53]) );
  CAN2X1 U7505 ( .A(\s10.addr[9] ), .B(n4167), .Z(\s10.SbusIn [60]) );
  CAN2XL U7506 ( .A(\s8.addr[17] ), .B(n4161), .Z(\s8.SbusIn [57]) );
  CAN2X1 U7507 ( .A(\s8.addr[15] ), .B(n4120), .Z(\s8.SbusIn [63]) );
  CAN2X1 U7508 ( .A(\s8.addr[15] ), .B(n3461), .Z(\s8.SbusIn [55]) );
  CAN2XL U7509 ( .A(\s8.addr[17] ), .B(n4157), .Z(\s8.addr [32]) );
  CAN2X1 U7510 ( .A(\s10.addr[9] ), .B(n4328), .Z(\s10.addr [25]) );
  CAN2XL U7511 ( .A(\s8.addr[17] ), .B(n4330), .Z(\s8.addr [2]) );
  CAN2X1 U7512 ( .A(\s8.addr[15] ), .B(n4201), .Z(\s8.addr [55]) );
  CAN2X1 U7513 ( .A(\s10.addr[9] ), .B(n4140), .Z(\s10.addr [63]) );
  CAN2X1 U7514 ( .A(\s8.addr[15] ), .B(n4160), .Z(\s8.addr [31]) );
  CAN2X1 U7515 ( .A(\s8.addr[15] ), .B(n4155), .Z(\s8.addr [49]) );
  CAN2X1 U7516 ( .A(\s8.addr[17] ), .B(n4165), .Z(\s8.addr [51]) );
  CAN2XL U7517 ( .A(\s8.addr[17] ), .B(n4131), .Z(\s8.addr [34]) );
  CAN2XL U7518 ( .A(\s8.en ), .B(n4176), .Z(\s8.addr [30]) );
  CAN2X1 U7519 ( .A(\s8.addr[17] ), .B(n3482), .Z(\s8.addr [60]) );
  CAN2XL U7520 ( .A(\s8.addr[17] ), .B(n4204), .Z(\s8.addr [38]) );
  CAN2XL U7521 ( .A(\s8.addr[17] ), .B(n3470), .Z(\s8.addr [44]) );
  CAN2XL U7522 ( .A(\s8.addr[17] ), .B(n3486), .Z(\s8.addr [40]) );
  CAN2XL U7523 ( .A(\s8.addr[17] ), .B(n3471), .Z(\s8.addr [41]) );
  CAN2X1 U7524 ( .A(\s7.addr[19] ), .B(n4196), .Z(\s7.SbusIn [37]) );
  CAN2XL U7525 ( .A(\s8.addr[17] ), .B(n4133), .Z(\s8.addr [28]) );
  CAN2XL U7526 ( .A(\s8.en ), .B(n4146), .Z(\s8.addr [47]) );
  CAN2XL U7527 ( .A(\s7.addr[16] ), .B(n4232), .Z(\s7.SbusIn [38]) );
  CAN2XL U7528 ( .A(\s7.addr[19] ), .B(n3475), .Z(\s7.addr [10]) );
  CAN2X1 U7529 ( .A(n4336), .B(n4175), .Z(\s7.SbusIn [54]) );
  CAN2X1 U7530 ( .A(\s7.addr[19] ), .B(n4174), .Z(\s7.addr [53]) );
  CAN2X1 U7531 ( .A(\s7.en ), .B(n4331), .Z(\s7.addr [20]) );
  CAN2XL U7532 ( .A(\s8.addr[15] ), .B(n4117), .Z(\s8.SbusIn [28]) );
  CAN2XL U7533 ( .A(\s8.addr[17] ), .B(n4159), .Z(\s8.SbusIn [56]) );
  CAN2XL U7534 ( .A(\s8.addr[17] ), .B(n3477), .Z(\s8.addr [59]) );
  CAN2XL U7535 ( .A(\s8.addr[17] ), .B(n4129), .Z(\s8.SbusIn [45]) );
  CAN2XL U7536 ( .A(\s6.addr [17]), .B(n4157), .Z(\s6.addr [32]) );
  CAN2XL U7537 ( .A(\s8.addr[17] ), .B(n4328), .Z(\s8.addr [25]) );
  CAN2XL U7538 ( .A(\s8.addr[17] ), .B(n4125), .Z(\s8.SbusIn [61]) );
  CAN2XL U7539 ( .A(\s1.addr [19]), .B(n3479), .Z(\s1.addr [62]) );
  CAN2XL U7540 ( .A(\s1.addr [19]), .B(n4175), .Z(\s1.SbusIn [54]) );
  CAN2XL U7541 ( .A(\s1.en ), .B(n4202), .Z(\s1.addr [58]) );
  CAN2XL U7542 ( .A(\s1.en ), .B(n3470), .Z(\s1.addr [44]) );
  CAN2XL U7543 ( .A(\s1.addr [19]), .B(n4148), .Z(\s1.addr [54]) );
  CAN2X1 U7544 ( .A(\s7.en ), .B(n4131), .Z(\s7.addr [34]) );
  CAN2X1 U7545 ( .A(\s7.en ), .B(n4124), .Z(\s7.addr [36]) );
  CAN2X1 U7546 ( .A(n4336), .B(n4136), .Z(\s7.addr [46]) );
  CAN2X1 U7547 ( .A(\s7.addr[16] ), .B(n4146), .Z(\s7.addr [47]) );
  CAN2XL U7548 ( .A(\s11.addr[17] ), .B(n3464), .Z(\s11.addr [37]) );
  CAN2XL U7549 ( .A(\s11.addr[19] ), .B(n4122), .Z(\s11.addr [43]) );
  CAN2XL U7550 ( .A(\s11.addr[19] ), .B(n4165), .Z(\s11.addr [51]) );
  CAN2XL U7551 ( .A(\s11.addr[17] ), .B(n4153), .Z(\s11.addr [42]) );
  CAN2XL U7552 ( .A(\s3.addr[14] ), .B(n4335), .Z(\s3.addr [8]) );
  CAN2XL U7553 ( .A(\s11.addr[19] ), .B(n4166), .Z(\s11.addr [52]) );
  CAN2XL U7554 ( .A(\s11.addr[19] ), .B(n3479), .Z(\s11.addr [62]) );
  CAN2XL U7555 ( .A(\s7.addr[16] ), .B(n4165), .Z(\s7.addr [51]) );
  CAN2XL U7556 ( .A(\s7.addr[19] ), .B(n4140), .Z(\s7.addr [63]) );
  CAN2XL U7557 ( .A(n4336), .B(n3470), .Z(\s7.addr [44]) );
  CAN2XL U7558 ( .A(\s7.en ), .B(n4166), .Z(\s7.addr [52]) );
  CNR2X1 U7559 ( .A(n4258), .B(n4326), .Z(\s13.addr [6]) );
  CAN2X1 U7560 ( .A(\s7.addr[16] ), .B(n4148), .Z(\s7.addr [54]) );
  CAN2X1 U7561 ( .A(\s7.en ), .B(n4133), .Z(\s7.addr [28]) );
  CAN2X1 U7562 ( .A(\s7.addr[19] ), .B(n4137), .Z(\s7.addr [48]) );
  CAN2X1 U7563 ( .A(\s14.addr [11]), .B(n4122), .Z(\s14.addr [43]) );
  CAN2X1 U7564 ( .A(\s9.addr[8] ), .B(n4195), .Z(\s9.addr [26]) );
  CAN2X1 U7565 ( .A(\s14.addr[18] ), .B(n4124), .Z(\s14.addr [36]) );
  CAN2X1 U7566 ( .A(\s14.addr[18] ), .B(n4146), .Z(\s14.addr [47]) );
  CAN2X1 U7567 ( .A(\s14.addr[18] ), .B(n4153), .Z(\s14.addr [42]) );
  CAN2X1 U7568 ( .A(\s14.addr[18] ), .B(n3470), .Z(\s14.addr [44]) );
  CAN2X1 U7569 ( .A(\s8.addr[17] ), .B(n4207), .Z(\s8.addr [57]) );
  CAN2XL U7570 ( .A(\s4.en ), .B(n4136), .Z(\s4.addr [46]) );
  CAN2XL U7571 ( .A(\s4.addr[14] ), .B(n4242), .Z(\s4.addr [56]) );
  CAN2XL U7572 ( .A(\s4.en ), .B(n4147), .Z(\s4.SbusIn [26]) );
  CAN2XL U7573 ( .A(\s4.addr[14] ), .B(n4161), .Z(\s4.SbusIn [57]) );
  CAN2XL U7574 ( .A(\s4.addr[14] ), .B(n4154), .Z(\s4.SbusIn [7]) );
  CAN2XL U7575 ( .A(\s4.addr[14] ), .B(n3487), .Z(\s4.SbusIn [16]) );
  CIVDX4 U7576 ( .A(n3457), .Z0(n3458), .Z1(n2740) );
  CIVX16 U7577 ( .A(n3458), .Z(n4256) );
  CNR2X1 U7578 ( .A(n4256), .B(n3459), .Z(\s2.addr [3]) );
  CAN2XL U7579 ( .A(n4405), .B(n3476), .Z(\s5.addr [5]) );
  CIVDX4 U7580 ( .A(n4188), .Z0(n4325), .Z1(\s0.addr [14]) );
  CNR2X1 U7581 ( .A(n4325), .B(n3459), .Z(\s0.addr [3]) );
  CAN2X1 U7582 ( .A(\s9.addr[16] ), .B(n4199), .Z(\s9.addr [24]) );
  CAN2XL U7583 ( .A(\s4.addr[14] ), .B(n4158), .Z(\s4.SbusIn [21]) );
  CAN2X1 U7584 ( .A(\s8.addr[15] ), .B(n4174), .Z(\s8.addr [53]) );
  CAN2XL U7585 ( .A(\s4.addr [19]), .B(n3476), .Z(\s4.addr [5]) );
  CAN2XL U7586 ( .A(\s4.addr[14] ), .B(n3486), .Z(\s4.addr [40]) );
  CAN2XL U7587 ( .A(\s4.addr[14] ), .B(n3462), .Z(\s4.addr [22]) );
  CAN2X1 U7588 ( .A(\s8.addr[15] ), .B(n4242), .Z(\s8.addr [56]) );
  CAN2X1 U7589 ( .A(\s8.addr[15] ), .B(n4134), .Z(\s8.addr [29]) );
  CAN2XL U7590 ( .A(\s4.addr[14] ), .B(n3460), .Z(\s4.SbusIn [27]) );
  CAN2X1 U7591 ( .A(\s3.addr[14] ), .B(n4154), .Z(\s3.SbusIn [7]) );
  CAN2XL U7592 ( .A(\s3.addr[14] ), .B(n3486), .Z(\s3.addr [40]) );
  CAN2XL U7593 ( .A(\s3.addr[9] ), .B(n4158), .Z(\s3.SbusIn [21]) );
  CAN2XL U7594 ( .A(\s4.en ), .B(n3469), .Z(\s4.SbusIn [5]) );
  CAN2XL U7595 ( .A(\s4.en ), .B(n4141), .Z(\s4.SbusIn [25]) );
  CAN2XL U7596 ( .A(\s6.en ), .B(n4131), .Z(\s6.addr [34]) );
  CIVDX4 U7597 ( .A(n4188), .Z0(n4327), .Z1(n4083) );
  CNR2X1 U7598 ( .A(n4327), .B(n4253), .Z(\s0.addr [5]) );
  CIVDX4 U7599 ( .A(n4188), .Z0(n4319), .Z1(\s0.addr[17] ) );
  CNR2X1 U7600 ( .A(n4319), .B(n3468), .Z(\s0.addr [1]) );
  CNR2X1 U7601 ( .A(n4317), .B(n4254), .Z(\s0.addr [4]) );
  CAN2XL U7602 ( .A(\s9.addr[7] ), .B(n4166), .Z(\s9.addr [52]) );
  CAN2XL U7603 ( .A(\s4.addr [19]), .B(n3470), .Z(\s4.addr [44]) );
  CAN2XL U7604 ( .A(\s4.addr [19]), .B(n4125), .Z(\s4.SbusIn [61]) );
  CAN2X1 U7605 ( .A(n4405), .B(n4179), .Z(\s5.addr [33]) );
  CAN2X1 U7606 ( .A(n1844), .B(n4153), .Z(\s5.addr [42]) );
  CAN2X1 U7607 ( .A(n5445), .B(n4207), .Z(\s5.addr [57]) );
  CAN2XL U7608 ( .A(\s1.addr[15] ), .B(n4140), .Z(\s1.addr [63]) );
  CAN2XL U7609 ( .A(\s1.addr[17] ), .B(n4200), .Z(\s1.SbusIn [3]) );
  CAN2XL U7610 ( .A(\s1.addr[17] ), .B(n4174), .Z(\s1.addr [53]) );
  CAN2XL U7611 ( .A(\s1.addr[17] ), .B(n4128), .Z(\s1.addr [21]) );
  CAN2XL U7612 ( .A(\s6.en ), .B(n4137), .Z(\s6.addr [48]) );
  CAN2XL U7613 ( .A(\s6.en ), .B(n3464), .Z(\s6.addr [37]) );
  CAN2XL U7614 ( .A(\s6.en ), .B(n3482), .Z(\s6.addr [60]) );
  CAN2XL U7615 ( .A(\s6.en ), .B(n4118), .Z(\s6.addr [23]) );
  CAN2XL U7616 ( .A(\s6.en ), .B(n4177), .Z(\s6.addr [39]) );
  CAN2XL U7617 ( .A(\s14.addr [11]), .B(n4119), .Z(\s14.SbusIn [31]) );
  CAN2XL U7618 ( .A(\s14.addr[17] ), .B(n4132), .Z(\s14.SbusIn [43]) );
  CAN2XL U7619 ( .A(\s14.addr [11]), .B(n4242), .Z(\s14.addr [56]) );
  CAN2XL U7620 ( .A(\s14.addr[17] ), .B(n4137), .Z(\s14.addr [48]) );
  CAN2XL U7621 ( .A(\s14.addr[17] ), .B(n4136), .Z(\s14.addr [46]) );
  CAN2XL U7622 ( .A(n4405), .B(n4242), .Z(\s5.addr [56]) );
  CAN2XL U7623 ( .A(n4405), .B(n3470), .Z(\s5.addr [44]) );
  CAN2XL U7624 ( .A(n4405), .B(n3460), .Z(\s5.SbusIn [27]) );
  CAN2XL U7625 ( .A(n1844), .B(n3486), .Z(\s5.addr [40]) );
  CAN2XL U7626 ( .A(\s6.en ), .B(n3480), .Z(\s6.SbusIn [49]) );
  CAN2XL U7627 ( .A(\s6.en ), .B(n4122), .Z(\s6.addr [43]) );
  CAN2XL U7628 ( .A(\s6.en ), .B(n4328), .Z(\s6.addr [25]) );
  CAN2XL U7629 ( .A(\s6.en ), .B(n4164), .Z(\s6.addr [50]) );
  CAN2XL U7630 ( .A(\s3.addr[9] ), .B(n4125), .Z(\s3.SbusIn [61]) );
  CAN2XL U7631 ( .A(\s3.addr[14] ), .B(n4119), .Z(\s3.SbusIn [31]) );
  CAN2XL U7632 ( .A(\s3.addr[14] ), .B(n4131), .Z(\s3.addr [34]) );
  CAN2XL U7633 ( .A(\s9.addr[8] ), .B(n4140), .Z(\s9.addr [63]) );
  CAN2XL U7634 ( .A(n4332), .B(n3486), .Z(\s11.addr [40]) );
  CAN2XL U7635 ( .A(\s12.addr[11] ), .B(n3485), .Z(\s12.addr [6]) );
  CAN2XL U7636 ( .A(\s4.addr [19]), .B(n4142), .Z(\s4.SbusIn [41]) );
  CAN2XL U7637 ( .A(\s4.addr[14] ), .B(n4131), .Z(\s4.addr [34]) );
  CAN2XL U7638 ( .A(\s4.addr[14] ), .B(n4151), .Z(\s4.addr [61]) );
  CAN2XL U7639 ( .A(\s4.en ), .B(n4215), .Z(\s4.SbusIn [36]) );
  CAN2XL U7640 ( .A(\s4.en ), .B(n4115), .Z(\s4.SbusIn [10]) );
  CAN2XL U7641 ( .A(\s4.en ), .B(n4130), .Z(\s4.SbusIn [59]) );
  CAN2XL U7642 ( .A(\s4.en ), .B(n4119), .Z(\s4.SbusIn [31]) );
  CAN2XL U7643 ( .A(\s4.addr[14] ), .B(n3479), .Z(\s4.addr [62]) );
  CAN2XL U7644 ( .A(\s4.en ), .B(n4156), .Z(\s4.SbusIn [33]) );
  CAN2XL U7645 ( .A(\s4.en ), .B(n3481), .Z(\s4.SbusIn [12]) );
  CAN2XL U7646 ( .A(\s4.en ), .B(n4152), .Z(\s4.SbusIn [19]) );
  CAN2XL U7647 ( .A(\s4.addr [19]), .B(n4168), .Z(\s4.SbusIn [58]) );
  CAN2XL U7648 ( .A(\s4.en ), .B(n4144), .Z(\s4.SbusIn [42]) );
  CAN2XL U7649 ( .A(\s4.en ), .B(n4165), .Z(\s4.addr [51]) );
  CAN2XL U7650 ( .A(\s4.en ), .B(n3480), .Z(\s4.SbusIn [49]) );
  CAN2XL U7651 ( .A(\s4.en ), .B(n4117), .Z(\s4.SbusIn [28]) );
  CAN2XL U7652 ( .A(\s4.en ), .B(n4126), .Z(\s4.SbusIn [62]) );
  CAN2XL U7653 ( .A(\s4.en ), .B(n4172), .Z(\s4.SbusIn [17]) );
  CAN2XL U7654 ( .A(\s4.en ), .B(n3474), .Z(\s4.SbusIn [14]) );
  CAN2XL U7655 ( .A(\s4.en ), .B(n3482), .Z(\s4.addr [60]) );
  CAN2XL U7656 ( .A(\s4.addr [19]), .B(n4175), .Z(\s4.SbusIn [54]) );
  CAN2XL U7657 ( .A(\s4.addr [19]), .B(n4170), .Z(\s4.SbusIn [53]) );
  CAN2XL U7658 ( .A(\s4.addr [19]), .B(n4193), .Z(\s4.SbusIn [9]) );
  CAN2XL U7659 ( .A(\s4.addr [19]), .B(n4190), .Z(\s4.SbusIn [1]) );
  CAN2XL U7660 ( .A(\s4.addr [19]), .B(n4243), .Z(\s4.SbusIn [4]) );
  CAN2XL U7661 ( .A(\s4.en ), .B(n3471), .Z(\s4.addr [41]) );
  CAN2XL U7662 ( .A(\s4.addr[14] ), .B(n4150), .Z(\s4.SbusIn [20]) );
  CAN2XL U7663 ( .A(\s4.addr [19]), .B(n4143), .Z(\s4.SbusIn [40]) );
  CAN2XL U7664 ( .A(\s4.en ), .B(n4160), .Z(\s4.addr [31]) );
  CAN2XL U7665 ( .A(\s4.addr[14] ), .B(n4192), .Z(\s4.SbusIn [2]) );
  CAN2XL U7666 ( .A(\s4.en ), .B(n4200), .Z(\s4.SbusIn [3]) );
  CAN2XL U7667 ( .A(\s4.en ), .B(n4120), .Z(\s4.SbusIn [63]) );
  CAN2XL U7668 ( .A(\s4.addr [19]), .B(n4149), .Z(\s4.SbusIn [24]) );
  CAN2XL U7669 ( .A(\s4.addr [19]), .B(n3461), .Z(\s4.SbusIn [55]) );
  CAN2XL U7670 ( .A(\s4.addr[14] ), .B(n4159), .Z(\s4.SbusIn [56]) );
  CAN2XL U7671 ( .A(\s4.en ), .B(n4123), .Z(\s4.SbusIn [13]) );
  CAN2XL U7672 ( .A(\s4.en ), .B(n4155), .Z(\s4.addr [49]) );
  CAN2XL U7673 ( .A(\s4.en ), .B(n4180), .Z(\s4.SbusIn [18]) );
  CAN2XL U7674 ( .A(\s4.en ), .B(n4134), .Z(\s4.addr [29]) );
  CAN2XL U7675 ( .A(\s4.en ), .B(n4201), .Z(\s4.addr [55]) );
  CAN2XL U7676 ( .A(\s4.addr [19]), .B(n4329), .Z(\s4.SbusIn [6]) );
  CAN2XL U7677 ( .A(\s4.addr [19]), .B(n4139), .Z(\s4.SbusIn [47]) );
  CAN2XL U7678 ( .A(\s4.addr [19]), .B(n4121), .Z(\s4.SbusIn [48]) );
  CAN2XL U7679 ( .A(\s4.addr[14] ), .B(n4129), .Z(\s4.SbusIn [45]) );
  CAN2XL U7680 ( .A(\s1.addr [19]), .B(n4131), .Z(\s1.addr [34]) );
  CAN2XL U7681 ( .A(\s1.addr[15] ), .B(n4328), .Z(\s1.addr [25]) );
  CAN2XL U7682 ( .A(\s1.en ), .B(n4124), .Z(\s1.addr [36]) );
  CAN2XL U7683 ( .A(\s6.en ), .B(n3485), .Z(\s6.addr [6]) );
  CAN2XL U7684 ( .A(\s6.en ), .B(n4162), .Z(\s6.addr [45]) );
  CAN2XL U7685 ( .A(\s14.addr [11]), .B(n4163), .Z(\s14.SbusIn [51]) );
  CAN2XL U7686 ( .A(\s14.addr[17] ), .B(n3485), .Z(\s14.addr [6]) );
  CAN2XL U7687 ( .A(n5445), .B(n4167), .Z(\s5.SbusIn [60]) );
  CAN2XL U7688 ( .A(n4405), .B(n4173), .Z(\s5.addr [35]) );
  CAN2XL U7689 ( .A(n4405), .B(n4176), .Z(\s5.addr [30]) );
  CAN2XL U7690 ( .A(n4405), .B(n4155), .Z(\s5.addr [49]) );
  CAN2XL U7691 ( .A(n4405), .B(n3487), .Z(\s5.SbusIn [16]) );
  CAN2XL U7692 ( .A(n1844), .B(n4142), .Z(\s5.SbusIn [41]) );
  CAN2XL U7693 ( .A(n5445), .B(n4128), .Z(\s5.addr [21]) );
  CAN2XL U7694 ( .A(n4405), .B(n4124), .Z(\s5.addr [36]) );
  CAN2XL U7695 ( .A(n4405), .B(n3466), .Z(\s5.SbusIn [52]) );
  CAN2XL U7696 ( .A(n4405), .B(n4133), .Z(\s5.addr [28]) );
  CAN2XL U7697 ( .A(n4405), .B(n3482), .Z(\s5.addr [60]) );
  CAN2XL U7698 ( .A(n1844), .B(n4139), .Z(\s5.SbusIn [47]) );
  CAN2XL U7699 ( .A(n5445), .B(n4136), .Z(\s5.addr [46]) );
  CAN2XL U7700 ( .A(n4405), .B(n4129), .Z(\s5.SbusIn [45]) );
  CAN2XL U7701 ( .A(n4405), .B(n4172), .Z(\s5.SbusIn [17]) );
  CAN2XL U7702 ( .A(n4405), .B(n4143), .Z(\s5.SbusIn [40]) );
  CAN2XL U7703 ( .A(\s7.addr[16] ), .B(n4155), .Z(\s7.addr [49]) );
  CAN2XL U7704 ( .A(\s7.addr[19] ), .B(n4134), .Z(\s7.addr [29]) );
  CAN2XL U7705 ( .A(\s7.en ), .B(n4202), .Z(\s7.addr [58]) );
  CAN2XL U7706 ( .A(\s7.en ), .B(n4128), .Z(\s7.addr [21]) );
  CAN2XL U7707 ( .A(\s3.addr[14] ), .B(n3466), .Z(\s3.SbusIn [52]) );
  CAN2XL U7708 ( .A(\s14.addr[17] ), .B(n4201), .Z(\s14.addr [55]) );
  CAN2XL U7709 ( .A(n4332), .B(n4141), .Z(\s11.SbusIn [25]) );
  CAN2XL U7710 ( .A(\s7.addr[16] ), .B(n4162), .Z(\s7.addr [45]) );
  CAN2XL U7711 ( .A(\s7.addr[19] ), .B(n4157), .Z(\s7.addr [32]) );
  CAN2XL U7712 ( .A(\s7.en ), .B(n4199), .Z(\s7.addr [24]) );
  CAN2XL U7713 ( .A(\s3.addr[14] ), .B(n3462), .Z(\s3.addr [22]) );
  CAN2XL U7714 ( .A(\s3.addr[14] ), .B(n4177), .Z(\s3.addr [39]) );
  CAN2XL U7715 ( .A(\s3.addr[14] ), .B(n4145), .Z(\s3.SbusIn [30]) );
  CAN2XL U7716 ( .A(\s3.addr[14] ), .B(n4164), .Z(\s3.addr [50]) );
  CAN2XL U7717 ( .A(\s3.addr[9] ), .B(n4197), .Z(\s3.SbusIn [29]) );
  CAN2XL U7718 ( .A(\s11.addr[19] ), .B(n3480), .Z(\s11.SbusIn [49]) );
  CAN2XL U7719 ( .A(\s3.addr [18]), .B(n4118), .Z(\s3.addr [23]) );
  CAN2XL U7720 ( .A(\s3.addr[14] ), .B(n4161), .Z(\s3.SbusIn [57]) );
  CAN2XL U7721 ( .A(n3463), .B(n3485), .Z(\s9.addr [6]) );
  CAN2XL U7722 ( .A(\s11.en ), .B(n3471), .Z(\s11.addr [41]) );
  CAN2XL U7723 ( .A(\s11.en ), .B(n4201), .Z(\s11.addr [55]) );
  CAN2XL U7724 ( .A(\s11.en ), .B(n4242), .Z(\s11.addr [56]) );
  CAN2XL U7725 ( .A(\s11.en ), .B(n4131), .Z(\s11.addr [34]) );
  CAN2XL U7726 ( .A(\s4.addr [19]), .B(n4137), .Z(\s4.addr [48]) );
  CAN2XL U7727 ( .A(\s4.addr[14] ), .B(n3464), .Z(\s4.addr [37]) );
  CAN2XL U7728 ( .A(\s4.addr[14] ), .B(n3472), .Z(\s4.SbusIn [46]) );
  CAN2XL U7729 ( .A(\s4.en ), .B(n4195), .Z(\s4.addr [26]) );
  CAN2XL U7730 ( .A(\s4.addr [19]), .B(n4328), .Z(\s4.addr [25]) );
  CAN2XL U7731 ( .A(\s4.en ), .B(n4133), .Z(\s4.addr [28]) );
  CAN2XL U7732 ( .A(\s4.en ), .B(n3477), .Z(\s4.addr [59]) );
  CAN2XL U7733 ( .A(\s4.en ), .B(n4185), .Z(\s4.SbusIn [0]) );
  CAN2XL U7734 ( .A(\s4.en ), .B(n4122), .Z(\s4.addr [43]) );
  CAN2XL U7735 ( .A(\s4.addr [19]), .B(n4138), .Z(\s4.SbusIn [44]) );
  CAN2XL U7736 ( .A(\s8.addr[17] ), .B(n4199), .Z(\s8.addr [24]) );
  CAN2XL U7737 ( .A(\s8.addr[17] ), .B(n4140), .Z(\s8.addr [63]) );
  CAN2XL U7738 ( .A(\s4.addr [19]), .B(n4169), .Z(\s4.SbusIn [15]) );
  CAN2XL U7739 ( .A(\s4.en ), .B(n3465), .Z(\s4.SbusIn [11]) );
  CAN2XL U7740 ( .A(\s4.addr [19]), .B(n4171), .Z(\s4.SbusIn [32]) );
  CAN2XL U7741 ( .A(\s4.addr [19]), .B(n4146), .Z(\s4.addr [47]) );
  CAN2XL U7742 ( .A(\s4.addr [19]), .B(n4179), .Z(\s4.addr [33]) );
  CAN2XL U7743 ( .A(\s4.addr[14] ), .B(n4118), .Z(\s4.addr [23]) );
  CAN2XL U7744 ( .A(\s4.addr[14] ), .B(n4331), .Z(\s4.addr [20]) );
  CAN2XL U7745 ( .A(\s4.en ), .B(n4127), .Z(\s4.SbusIn [50]) );
  CAN2XL U7746 ( .A(\s8.addr[17] ), .B(n4162), .Z(\s8.addr [45]) );
  CAN2XL U7747 ( .A(\s4.addr [19]), .B(n4232), .Z(\s4.SbusIn [38]) );
  CAN2XL U7748 ( .A(\s4.addr [19]), .B(n4167), .Z(\s4.SbusIn [60]) );
  CAN2XL U7749 ( .A(\s4.addr[14] ), .B(n4128), .Z(\s4.addr [21]) );
  CAN2XL U7750 ( .A(\s4.addr[14] ), .B(n4176), .Z(\s4.addr [30]) );
  CAN2XL U7751 ( .A(\s4.addr [19]), .B(n4174), .Z(\s4.addr [53]) );
  CAN2XL U7752 ( .A(\s4.en ), .B(n4173), .Z(\s4.addr [35]) );
  CAN2XL U7753 ( .A(\s4.en ), .B(n4196), .Z(\s4.SbusIn [37]) );
  CAN2XL U7754 ( .A(\s4.addr [19]), .B(n4177), .Z(\s4.addr [39]) );
  CAN2XL U7755 ( .A(\s4.addr[14] ), .B(n4157), .Z(\s4.addr [32]) );
  CAN2XL U7756 ( .A(\s4.addr[14] ), .B(n4163), .Z(\s4.SbusIn [51]) );
  CAN2XL U7757 ( .A(\s4.addr [19]), .B(n4145), .Z(\s4.SbusIn [30]) );
  CAN2XL U7758 ( .A(\s4.addr[14] ), .B(n3473), .Z(\s4.SbusIn [22]) );
  CAN2XL U7759 ( .A(\s4.addr[14] ), .B(n4140), .Z(\s4.addr [63]) );
  CAN2XL U7760 ( .A(\s4.addr[14] ), .B(n3467), .Z(\s4.addr [27]) );
  CAN2XL U7761 ( .A(\s4.en ), .B(n4148), .Z(\s4.addr [54]) );
  CAN2XL U7762 ( .A(\s4.en ), .B(n4202), .Z(\s4.addr [58]) );
  CAN2XL U7763 ( .A(\s4.addr[14] ), .B(n4124), .Z(\s4.addr [36]) );
  CAN2XL U7764 ( .A(\s4.addr [19]), .B(n4132), .Z(\s4.SbusIn [43]) );
  CAN2XL U7765 ( .A(\s4.addr[14] ), .B(n4135), .Z(\s4.SbusIn [39]) );
  CAN2XL U7766 ( .A(\s4.en ), .B(n4153), .Z(\s4.addr [42]) );
  CAN2XL U7767 ( .A(\s4.addr [19]), .B(n4199), .Z(\s4.addr [24]) );
  CAN2XL U7768 ( .A(\s4.addr[14] ), .B(n3466), .Z(\s4.SbusIn [52]) );
  CAN2XL U7769 ( .A(\s4.en ), .B(n4207), .Z(\s4.addr [57]) );
  CAN2XL U7770 ( .A(\s4.en ), .B(n4178), .Z(\s4.SbusIn [34]) );
  CAN2XL U7771 ( .A(\s4.addr [19]), .B(n4162), .Z(\s4.addr [45]) );
  CAN2XL U7772 ( .A(\s4.en ), .B(n4116), .Z(\s4.SbusIn [8]) );
  CAN2XL U7773 ( .A(\s4.en ), .B(n4197), .Z(\s4.SbusIn [29]) );
  CAN2XL U7774 ( .A(\s4.addr [19]), .B(n3483), .Z(\s4.SbusIn [23]) );
  CAN2XL U7775 ( .A(\s4.addr [19]), .B(n4166), .Z(\s4.addr [52]) );
  CAN2XL U7776 ( .A(\s4.addr[14] ), .B(n4164), .Z(\s4.addr [50]) );
  CAN2XL U7777 ( .A(\s4.en ), .B(n4204), .Z(\s4.addr [38]) );
  CAN2XL U7778 ( .A(\s1.addr[17] ), .B(n4177), .Z(\s1.addr [39]) );
  CAN2XL U7779 ( .A(\s1.en ), .B(n4171), .Z(\s1.SbusIn [32]) );
  CAN2XL U7780 ( .A(\s1.en ), .B(n4204), .Z(\s1.addr [38]) );
  CAN2XL U7781 ( .A(\s1.addr[15] ), .B(n4138), .Z(\s1.SbusIn [44]) );
  CAN2XL U7782 ( .A(\s1.addr[17] ), .B(n4195), .Z(\s1.addr [26]) );
  CAN2XL U7783 ( .A(\s1.addr[15] ), .B(n3467), .Z(\s1.addr [27]) );
  CAN2XL U7784 ( .A(\s1.addr[17] ), .B(n4173), .Z(\s1.addr [35]) );
  CNR2X1 U7785 ( .A(n4256), .B(n3468), .Z(\s2.addr [1]) );
  CAN2XL U7786 ( .A(\s3.addr[14] ), .B(n3469), .Z(\s3.SbusIn [5]) );
  CAN2XL U7787 ( .A(\s3.addr[9] ), .B(n3480), .Z(\s3.SbusIn [49]) );
  CAN2XL U7788 ( .A(\s3.addr[14] ), .B(n4242), .Z(\s3.addr [56]) );
  CAN2XL U7789 ( .A(\s3.addr [18]), .B(n4201), .Z(\s3.addr [55]) );
  CAN2XL U7790 ( .A(\s3.addr[14] ), .B(n4155), .Z(\s3.addr [49]) );
  CAN2XL U7791 ( .A(\s3.addr[14] ), .B(n4129), .Z(\s3.SbusIn [45]) );
  CAN2XL U7792 ( .A(\s3.addr [18]), .B(n3470), .Z(\s3.addr [44]) );
  CAN2XL U7793 ( .A(n1844), .B(n4157), .Z(\s5.addr [32]) );
  CAN2XL U7794 ( .A(n5445), .B(n4195), .Z(\s5.addr [26]) );
  CAN2XL U7795 ( .A(n4405), .B(n3473), .Z(\s5.SbusIn [22]) );
  CAN2XL U7796 ( .A(n4405), .B(n4237), .Z(\s5.SbusIn [35]) );
  CAN2XL U7797 ( .A(\s3.addr[9] ), .B(n3471), .Z(\s3.addr [41]) );
  CAN2XL U7798 ( .A(\s3.addr [18]), .B(n4328), .Z(\s3.addr [25]) );
  CAN2XL U7799 ( .A(\s3.addr [18]), .B(n4150), .Z(\s3.SbusIn [20]) );
  CAN2XL U7800 ( .A(\s3.addr[9] ), .B(n3472), .Z(\s3.SbusIn [46]) );
  CAN2XL U7801 ( .A(\s3.addr[9] ), .B(n4170), .Z(\s3.SbusIn [53]) );
  CAN2XL U7802 ( .A(\s3.addr[9] ), .B(n4163), .Z(\s3.SbusIn [51]) );
  CAN2XL U7803 ( .A(\s3.addr[9] ), .B(n4172), .Z(\s3.SbusIn [17]) );
  CAN2XL U7804 ( .A(\s3.addr [18]), .B(n4135), .Z(\s3.SbusIn [39]) );
  CAN2XL U7805 ( .A(\s3.addr[14] ), .B(n4149), .Z(\s3.SbusIn [24]) );
  CAN2XL U7806 ( .A(\s3.addr[14] ), .B(n4144), .Z(\s3.SbusIn [42]) );
  CAN2XL U7807 ( .A(\s3.addr[9] ), .B(n4151), .Z(\s3.addr [61]) );
  CAN2XL U7808 ( .A(\s14.addr[17] ), .B(n4162), .Z(\s14.addr [45]) );
  CAN2XL U7809 ( .A(n4332), .B(n3476), .Z(\s11.addr [5]) );
  CAN2XL U7810 ( .A(n4332), .B(n4176), .Z(\s11.addr [30]) );
  CAN2XL U7811 ( .A(n4332), .B(n4178), .Z(\s11.SbusIn [34]) );
  CAN2XL U7812 ( .A(n4332), .B(n4177), .Z(\s11.addr [39]) );
  CAN2XL U7813 ( .A(n4332), .B(n3473), .Z(\s11.SbusIn [22]) );
  CAN2XL U7814 ( .A(n4332), .B(n4193), .Z(\s11.SbusIn [9]) );
  CAN2XL U7815 ( .A(n4332), .B(n3477), .Z(\s11.addr [59]) );
  CAN2XL U7816 ( .A(n4332), .B(n4185), .Z(\s11.SbusIn [0]) );
  CAN2XL U7817 ( .A(n4332), .B(n4162), .Z(\s11.addr [45]) );
  CAN2XL U7818 ( .A(n4332), .B(n4127), .Z(\s11.SbusIn [50]) );
  CAN2XL U7819 ( .A(\s3.addr[14] ), .B(n4196), .Z(\s3.SbusIn [37]) );
  CAN2XL U7820 ( .A(\s3.addr[9] ), .B(n4152), .Z(\s3.SbusIn [19]) );
  CAN2XL U7821 ( .A(\s3.addr [18]), .B(n3474), .Z(\s3.SbusIn [14]) );
  CAN2XL U7822 ( .A(\s3.addr[14] ), .B(n4178), .Z(\s3.SbusIn [34]) );
  CAN2XL U7823 ( .A(\s11.addr[19] ), .B(n3475), .Z(\s11.addr [10]) );
  CAN2XL U7824 ( .A(\s7.addr[19] ), .B(n4195), .Z(\s7.addr [26]) );
  CAN2XL U7825 ( .A(\s3.addr[9] ), .B(n3476), .Z(\s3.addr [5]) );
  CAN2XL U7826 ( .A(\s11.en ), .B(n4133), .Z(\s11.addr [28]) );
  CAN2XL U7827 ( .A(\s11.en ), .B(n4151), .Z(\s11.addr [61]) );
  CAN2XL U7828 ( .A(\s11.en ), .B(n4157), .Z(\s11.addr [32]) );
  CAN2XL U7829 ( .A(\s11.en ), .B(n4202), .Z(\s11.addr [58]) );
  CAN2XL U7830 ( .A(\s11.en ), .B(n4207), .Z(\s11.addr [57]) );
  CAN2XL U7831 ( .A(\s3.addr[9] ), .B(n4136), .Z(\s3.addr [46]) );
  CAN2XL U7832 ( .A(\s3.addr[14] ), .B(n4185), .Z(\s3.SbusIn [0]) );
  CAN2XL U7833 ( .A(\s3.addr[14] ), .B(n4171), .Z(\s3.SbusIn [32]) );
  CAN2XL U7834 ( .A(\s3.addr[14] ), .B(n4199), .Z(\s3.addr [24]) );
  CAN2XL U7835 ( .A(\s10.en ), .B(n3477), .Z(\s10.addr [59]) );
  CAN2XL U7836 ( .A(\s10.en ), .B(n4331), .Z(\s10.addr [20]) );
  CAN2XL U7837 ( .A(\s10.en ), .B(n4174), .Z(\s10.addr [53]) );
  CAN2XL U7838 ( .A(\s10.en ), .B(n4118), .Z(\s10.addr [23]) );
  CAN2XL U7839 ( .A(\s10.en ), .B(n4148), .Z(\s10.addr [54]) );
  CAN2XL U7840 ( .A(\s11.en ), .B(n4179), .Z(\s11.addr [33]) );
  CAN2XL U7841 ( .A(n4332), .B(n3487), .Z(\s11.SbusIn [16]) );
  CAN2XL U7842 ( .A(n4332), .B(n4164), .Z(\s11.addr [50]) );
  CAN2XL U7843 ( .A(n4332), .B(n4146), .Z(\s11.addr [47]) );
  CAN2XL U7844 ( .A(n4332), .B(n4174), .Z(\s11.addr [53]) );
  CAN2XL U7845 ( .A(n4332), .B(n4204), .Z(\s11.addr [38]) );
  CAN2XL U7846 ( .A(n4332), .B(n4148), .Z(\s11.addr [54]) );
  CAN2XL U7847 ( .A(\s11.en ), .B(n4140), .Z(\s11.addr [63]) );
  CAN2XL U7848 ( .A(n4332), .B(n4147), .Z(\s11.SbusIn [26]) );
  CAN2XL U7849 ( .A(\s8.addr[15] ), .B(n3478), .Z(\s8.addr [6]) );
  CAN2XL U7850 ( .A(\s7.addr[16] ), .B(n4330), .Z(\s7.addr [2]) );
  CAN2XL U7851 ( .A(\s10.addr [17]), .B(n4164), .Z(\s10.addr [50]) );
  CAN2XL U7852 ( .A(\s3.addr[14] ), .B(n3487), .Z(\s3.SbusIn [16]) );
  CAN2XL U7853 ( .A(\s3.addr[9] ), .B(n4147), .Z(\s3.SbusIn [26]) );
  CAN2XL U7854 ( .A(\s3.addr [18]), .B(n4141), .Z(\s3.SbusIn [25]) );
  CAN2XL U7855 ( .A(\s3.addr[14] ), .B(n4159), .Z(\s3.SbusIn [56]) );
  CAN2XL U7856 ( .A(\s3.addr[14] ), .B(n4232), .Z(\s3.SbusIn [38]) );
  CAN2XL U7857 ( .A(\s3.addr [18]), .B(n3479), .Z(\s3.addr [62]) );
  CAN2XL U7858 ( .A(n4405), .B(n4146), .Z(\s5.addr [47]) );
  CAN2XL U7859 ( .A(n4405), .B(n3480), .Z(\s5.SbusIn [49]) );
  CAN2XL U7860 ( .A(n1844), .B(n4196), .Z(\s5.SbusIn [37]) );
  CAN2XL U7861 ( .A(n5445), .B(n4190), .Z(\s5.SbusIn [1]) );
  CAN2XL U7862 ( .A(n4405), .B(n4152), .Z(\s5.SbusIn [19]) );
  CAN2XL U7863 ( .A(n4405), .B(n4123), .Z(\s5.SbusIn [13]) );
  CAN2XL U7864 ( .A(n4405), .B(n3481), .Z(\s5.SbusIn [12]) );
  CAN2XL U7865 ( .A(n4405), .B(n4178), .Z(\s5.SbusIn [34]) );
  CAN2XL U7866 ( .A(n1844), .B(n4201), .Z(\s5.addr [55]) );
  CAN2XL U7867 ( .A(n5445), .B(n4116), .Z(\s5.SbusIn [8]) );
  CAN2XL U7868 ( .A(n4405), .B(n4162), .Z(\s5.addr [45]) );
  CAN2XL U7869 ( .A(\s3.addr[9] ), .B(n4179), .Z(\s3.addr [33]) );
  CAN2XL U7870 ( .A(\s3.addr[14] ), .B(n4207), .Z(\s3.addr [57]) );
  CAN2XL U7871 ( .A(\s6.addr [17]), .B(n4330), .Z(\s6.addr [2]) );
  CAN2XL U7872 ( .A(\s3.addr[14] ), .B(n4176), .Z(\s3.addr [30]) );
  CAN2XL U7873 ( .A(\s3.addr[14] ), .B(n4202), .Z(\s3.addr [58]) );
  CAN2XL U7874 ( .A(\s3.addr [18]), .B(n4190), .Z(\s3.SbusIn [1]) );
  CAN2XL U7875 ( .A(\s3.addr[14] ), .B(n4134), .Z(\s3.addr [29]) );
  CAN2XL U7876 ( .A(\s3.addr[14] ), .B(n4142), .Z(\s3.SbusIn [41]) );
  CAN2XL U7877 ( .A(\s3.addr [18]), .B(n3482), .Z(\s3.addr [60]) );
  CAN2XL U7878 ( .A(\s3.addr[9] ), .B(n4192), .Z(\s3.SbusIn [2]) );
  CAN2XL U7879 ( .A(\s3.addr[14] ), .B(n4127), .Z(\s3.SbusIn [50]) );
  CAN2XL U7880 ( .A(\s3.addr[14] ), .B(n4128), .Z(\s3.addr [21]) );
  CAN2XL U7881 ( .A(\s3.addr[14] ), .B(n4204), .Z(\s3.addr [38]) );
  CAN2XL U7882 ( .A(\s3.addr[14] ), .B(n4195), .Z(\s3.addr [26]) );
  CAN2XL U7883 ( .A(\s3.addr[14] ), .B(n4117), .Z(\s3.SbusIn [28]) );
  CAN2XL U7884 ( .A(\s3.addr[14] ), .B(n4132), .Z(\s3.SbusIn [43]) );
  CAN2XL U7885 ( .A(\s3.addr[14] ), .B(n3483), .Z(\s3.SbusIn [23]) );
  CAN2XL U7886 ( .A(\s3.addr [18]), .B(n4160), .Z(\s3.addr [31]) );
  CAN2XL U7887 ( .A(\s3.addr[14] ), .B(n3485), .Z(\s3.addr [6]) );
  CAN2XL U7888 ( .A(\s3.addr[14] ), .B(n4180), .Z(\s3.SbusIn [18]) );
  CAN2XL U7889 ( .A(\s3.addr[14] ), .B(n4139), .Z(\s3.SbusIn [47]) );
  CAN2XL U7890 ( .A(\s3.addr[14] ), .B(n4124), .Z(\s3.addr [36]) );
  CAN2XL U7891 ( .A(\s11.addr[17] ), .B(n3484), .Z(\s11.addr [11]) );
  CAN2XL U7892 ( .A(\s11.en ), .B(n3485), .Z(\s11.addr [6]) );
  CAN2XL U7893 ( .A(\s10.en ), .B(n4195), .Z(\s10.addr [26]) );
  CAN2XL U7894 ( .A(\s11.en ), .B(n4330), .Z(\s11.addr [2]) );
  CAN2XL U7895 ( .A(\s10.addr[9] ), .B(n4131), .Z(\s10.addr [34]) );
  CAN2XL U7896 ( .A(\s10.addr[9] ), .B(n4136), .Z(\s10.addr [46]) );
  CAN2XL U7897 ( .A(\s10.en ), .B(n3486), .Z(\s10.addr [40]) );
  CAN2XL U7898 ( .A(\s10.en ), .B(n4242), .Z(\s10.addr [56]) );
  CAN2XL U7899 ( .A(\s10.en ), .B(n4165), .Z(\s10.addr [51]) );
  CAN2XL U7900 ( .A(\s10.en ), .B(n4146), .Z(\s10.addr [47]) );
  CAN2XL U7901 ( .A(\s10.en ), .B(n4202), .Z(\s10.addr [58]) );
  CAN2XL U7902 ( .A(\s10.en ), .B(n4137), .Z(\s10.addr [48]) );
  CAN2XL U7903 ( .A(\s10.en ), .B(n4162), .Z(\s10.addr [45]) );
  CAN2XL U7904 ( .A(\s10.en ), .B(n4176), .Z(\s10.addr [30]) );
  CAN2XL U7905 ( .A(\s10.en ), .B(n4151), .Z(\s10.addr [61]) );
  CAN2XL U7906 ( .A(\s10.en ), .B(n4330), .Z(\s10.addr [2]) );
  CAN2XL U7907 ( .A(\s10.en ), .B(n4204), .Z(\s10.addr [38]) );
  CAN2XL U7908 ( .A(n4405), .B(n4330), .Z(\s5.addr [2]) );
  CAN2X1 U7909 ( .A(\s9.addr[7] ), .B(n4202), .Z(\s9.addr [58]) );
  CAN2X1 U7910 ( .A(n5590), .B(n4128), .Z(\s9.addr [21]) );
  CAN2XL U7911 ( .A(\s14.addr[18] ), .B(n4335), .Z(\s14.addr [8]) );
  CAN2XL U7912 ( .A(\s12.addr[11] ), .B(n4335), .Z(\s12.addr [8]) );
  CAN2X1 U7913 ( .A(\s8.addr[15] ), .B(n3487), .Z(\s8.SbusIn [16]) );
  CAN2X1 U7914 ( .A(\s7.addr[19] ), .B(n3487), .Z(\s7.SbusIn [16]) );
  CAOR2XL U7915 ( .A(\s1.addr [19]), .B(\s1.dbus_out [15]), .C(n4072), .D(
        \s7.dbus_out [15]), .Z(n3489) );
  CAOR2XL U7916 ( .A(\c1.Breset ), .B(data_stm_d[15]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [15]), .Z(n3488) );
  CANR3XL U7917 ( .A(\s6.en ), .B(\s6.dbus_out [15]), .C(n3489), .D(n3488), 
        .Z(n3498) );
  CND2X1 U7918 ( .A(n4098), .B(\s10.dbus_out [15]), .Z(n3493) );
  CANR2XL U7919 ( .A(n4078), .B(\s5.dbus_out [15]), .C(n4091), .D(
        \s4.dbus_out [15]), .Z(n3492) );
  CANR2XL U7920 ( .A(\s14.dbus_out [15]), .B(\s14.addr [11]), .C(
        \s12.dbus_out [15]), .D(n1840), .Z(n3491) );
  CND2XL U7921 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [15]), .Z(n3490) );
  CAN4X1 U7922 ( .A(n3493), .B(n3492), .C(n3491), .D(n3490), .Z(n3497) );
  CAOR2XL U7923 ( .A(\s9.dbus_out [15]), .B(\s9.addr[7] ), .C(n4083), .D(
        \s0.dbus_out [15]), .Z(n3494) );
  CANR1XL U7924 ( .A(n4108), .B(\s11.dbus_out [15]), .C(n3494), .Z(n3496) );
  CANR2X1 U7925 ( .A(n4110), .B(\s13.dbus_out [15]), .C(n4085), .D(
        \s8.dbus_out [15]), .Z(n3495) );
  CND4X1 U7926 ( .A(n3498), .B(n3497), .C(n3496), .D(n3495), .Z(n1739) );
  CAOR2X1 U7927 ( .A(n4095), .B(\s1.dbus_out [1]), .C(n4072), .D(
        \s7.dbus_out [1]), .Z(n3500) );
  CAOR2XL U7928 ( .A(\c1.Breset ), .B(data_stm_d[1]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [1]), .Z(n3499) );
  CANR3X1 U7929 ( .A(\s6.addr [17]), .B(\s6.dbus_out [1]), .C(n3500), .D(n3499), .Z(n3509) );
  CND2X1 U7930 ( .A(n4098), .B(\s10.dbus_out [1]), .Z(n3504) );
  CNIVX2 U7931 ( .A(\s5.addr[14] ), .Z(n4078) );
  CANR2X1 U7932 ( .A(n4078), .B(\s5.dbus_out [1]), .C(n4091), .D(
        \s4.dbus_out [1]), .Z(n3503) );
  CANR2X1 U7933 ( .A(n4092), .B(\s14.dbus_out [1]), .C(\s12.dbus_out [1]), .D(
        n4099), .Z(n3502) );
  CND2XL U7934 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [1]), .Z(n3501) );
  CAN4X1 U7935 ( .A(n3504), .B(n3503), .C(n3502), .D(n3501), .Z(n3508) );
  CAOR2XL U7936 ( .A(\s9.dbus_out [1]), .B(\s9.addr[16] ), .C(n3975), .D(
        \s0.dbus_out [1]), .Z(n3505) );
  CANR1XL U7937 ( .A(\s11.dbus_out [1]), .B(\s11.addr[17] ), .C(n3505), .Z(
        n3507) );
  CANR2X1 U7938 ( .A(n4110), .B(\s13.dbus_out [1]), .C(n4085), .D(
        \s8.dbus_out [1]), .Z(n3506) );
  CND4X1 U7939 ( .A(n3509), .B(n3508), .C(n3507), .D(n3506), .Z(n1753) );
  CAOR2XL U7940 ( .A(n4090), .B(\s1.dbus_out [36]), .C(n4094), .D(
        \s7.dbus_out [36]), .Z(n3511) );
  CAOR2XL U7941 ( .A(\c1.Breset ), .B(data_stm_d[36]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [36]), .Z(n3510) );
  CANR3X1 U7942 ( .A(\s6.addr [17]), .B(\s6.dbus_out [36]), .C(n3511), .D(
        n3510), .Z(n3521) );
  CNR2IX1 U7943 ( .B(\s10.dbus_out [36]), .A(n4076), .Z(n3512) );
  CIVX2 U7944 ( .A(n3512), .Z(n3516) );
  CANR2XL U7945 ( .A(n4078), .B(\s5.dbus_out [36]), .C(n4077), .D(
        \s4.dbus_out [36]), .Z(n3515) );
  CANR2X1 U7946 ( .A(n4100), .B(\s14.dbus_out [36]), .C(\s12.dbus_out [36]), 
        .D(n4099), .Z(n3514) );
  CND2XL U7947 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [36]), .Z(n3513) );
  CAN4X1 U7948 ( .A(n3516), .B(n3515), .C(n3514), .D(n3513), .Z(n3520) );
  CAOR2XL U7949 ( .A(\s9.dbus_out [36]), .B(\s9.en ), .C(\s0.addr [12]), .D(
        \s0.dbus_out [36]), .Z(n3517) );
  CANR1XL U7950 ( .A(n4093), .B(\s11.dbus_out [36]), .C(n3517), .Z(n3519) );
  CANR2XL U7951 ( .A(n4110), .B(\s13.dbus_out [36]), .C(n4085), .D(
        \s8.dbus_out [36]), .Z(n3518) );
  CND4X1 U7952 ( .A(n3521), .B(n3520), .C(n3519), .D(n3518), .Z(n1718) );
  CNIVX1 U7953 ( .A(n1843), .Z(n4016) );
  CIVDX4 U7954 ( .A(n4188), .Z0(n4317), .Z1(n3963) );
  CAOR2XL U7955 ( .A(n4090), .B(\s1.dbus_out [61]), .C(n4094), .D(
        \s7.dbus_out [61]), .Z(n3523) );
  CAOR2XL U7956 ( .A(\c1.Breset ), .B(data_stm_d[61]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [61]), .Z(n3522) );
  CANR3X1 U7957 ( .A(n4075), .B(\s6.dbus_out [61]), .C(n3523), .D(n3522), .Z(
        n3532) );
  CND2X1 U7958 ( .A(n4098), .B(\s10.dbus_out [61]), .Z(n3527) );
  CANR2XL U7959 ( .A(n4078), .B(\s5.dbus_out [61]), .C(n4091), .D(
        \s4.dbus_out [61]), .Z(n3526) );
  CANR2XL U7960 ( .A(\s14.dbus_out [61]), .B(\s14.addr[16] ), .C(
        \s12.dbus_out [61]), .D(n4099), .Z(n3525) );
  CND2X1 U7961 ( .A(n4101), .B(\s3.dbus_out [61]), .Z(n3524) );
  CAN4X1 U7962 ( .A(n3527), .B(n3526), .C(n3525), .D(n3524), .Z(n3531) );
  CNIVX1 U7963 ( .A(\s11.addr[17] ), .Z(n3872) );
  CAOR2XL U7964 ( .A(\s9.dbus_out [61]), .B(\s9.addr[16] ), .C(n3940), .D(
        \s0.dbus_out [61]), .Z(n3528) );
  CANR1XL U7965 ( .A(\s11.dbus_out [61]), .B(n3872), .C(n3528), .Z(n3530) );
  CANR2XL U7966 ( .A(n4110), .B(\s13.dbus_out [61]), .C(n4109), .D(
        \s8.dbus_out [61]), .Z(n3529) );
  CND4X1 U7967 ( .A(n3532), .B(n3531), .C(n3530), .D(n3529), .Z(n1693) );
  CAOR2X1 U7968 ( .A(n4090), .B(\s1.dbus_out [35]), .C(n4072), .D(
        \s7.dbus_out [35]), .Z(n3534) );
  CAOR2XL U7969 ( .A(\c1.Breset ), .B(data_stm_d[35]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [35]), .Z(n3533) );
  CANR3XL U7970 ( .A(\s6.addr [17]), .B(\s6.dbus_out [35]), .C(n3534), .D(
        n3533), .Z(n3543) );
  CND2XL U7971 ( .A(n4098), .B(\s10.dbus_out [35]), .Z(n3538) );
  CANR2XL U7972 ( .A(n4078), .B(\s5.dbus_out [35]), .C(n4091), .D(
        \s4.dbus_out [35]), .Z(n3537) );
  CANR2XL U7973 ( .A(n4100), .B(\s14.dbus_out [35]), .C(\s12.dbus_out [35]), 
        .D(n1843), .Z(n3536) );
  CND2XL U7974 ( .A(n4101), .B(\s3.dbus_out [35]), .Z(n3535) );
  CAN4X1 U7975 ( .A(n3538), .B(n3537), .C(n3536), .D(n3535), .Z(n3542) );
  CAOR2XL U7976 ( .A(\s9.dbus_out [35]), .B(\s9.addr[8] ), .C(\s0.addr [12]), 
        .D(\s0.dbus_out [35]), .Z(n3539) );
  CANR1XL U7977 ( .A(n4108), .B(\s11.dbus_out [35]), .C(n3539), .Z(n3541) );
  CANR2X1 U7978 ( .A(n4110), .B(\s13.dbus_out [35]), .C(n4085), .D(
        \s8.dbus_out [35]), .Z(n3540) );
  CND4X1 U7979 ( .A(n3543), .B(n3542), .C(n3541), .D(n3540), .Z(n1719) );
  CAOR2XL U7980 ( .A(n4090), .B(\s1.dbus_out [48]), .C(n4072), .D(
        \s7.dbus_out [48]), .Z(n3545) );
  CAOR2XL U7981 ( .A(\c1.Breset ), .B(data_stm_d[48]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [48]), .Z(n3544) );
  CANR3XL U7982 ( .A(n4062), .B(\s6.dbus_out [48]), .C(n3545), .D(n3544), .Z(
        n3554) );
  CND2X1 U7983 ( .A(n4098), .B(\s10.dbus_out [48]), .Z(n3549) );
  CANR2XL U7984 ( .A(n4078), .B(\s5.dbus_out [48]), .C(\s4.addr [19]), .D(
        \s4.dbus_out [48]), .Z(n3548) );
  CANR2XL U7985 ( .A(\s14.addr[16] ), .B(\s14.dbus_out [48]), .C(
        \s12.dbus_out [48]), .D(n4099), .Z(n3547) );
  CND2XL U7986 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [48]), .Z(n3546) );
  CAN4X1 U7987 ( .A(n3549), .B(n3548), .C(n3547), .D(n3546), .Z(n3553) );
  CAOR2XL U7988 ( .A(\s9.dbus_out [48]), .B(\s9.addr[16] ), .C(n3963), .D(
        \s0.dbus_out [48]), .Z(n3550) );
  CANR1XL U7989 ( .A(n4093), .B(\s11.dbus_out [48]), .C(n3550), .Z(n3552) );
  CANR2X1 U7990 ( .A(n4110), .B(\s13.dbus_out [48]), .C(n4085), .D(
        \s8.dbus_out [48]), .Z(n3551) );
  CND4X1 U7991 ( .A(n3554), .B(n3553), .C(n3552), .D(n3551), .Z(n1706) );
  CAOR2XL U7992 ( .A(\s1.addr [19]), .B(\s1.dbus_out [47]), .C(n4094), .D(
        \s7.dbus_out [47]), .Z(n3556) );
  CAOR2XL U7993 ( .A(\c1.Breset ), .B(data_stm_d[47]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [47]), .Z(n3555) );
  CANR3XL U7994 ( .A(n4062), .B(\s6.dbus_out [47]), .C(n3556), .D(n3555), .Z(
        n3565) );
  CND2XL U7995 ( .A(n4098), .B(\s10.dbus_out [47]), .Z(n3560) );
  CANR2XL U7996 ( .A(n4078), .B(\s5.dbus_out [47]), .C(n4077), .D(
        \s4.dbus_out [47]), .Z(n3559) );
  CANR2X1 U7997 ( .A(n4100), .B(\s14.dbus_out [47]), .C(\s12.dbus_out [47]), 
        .D(n4099), .Z(n3558) );
  CND2X1 U7998 ( .A(n4101), .B(\s3.dbus_out [47]), .Z(n3557) );
  CAN4X1 U7999 ( .A(n3560), .B(n3559), .C(n3558), .D(n3557), .Z(n3564) );
  CAOR2XL U8000 ( .A(\s9.dbus_out [47]), .B(\s9.en ), .C(n4106), .D(
        \s0.dbus_out [47]), .Z(n3561) );
  CANR1XL U8001 ( .A(n4093), .B(\s11.dbus_out [47]), .C(n3561), .Z(n3563) );
  CANR2X1 U8002 ( .A(n4110), .B(\s13.dbus_out [47]), .C(n4085), .D(
        \s8.dbus_out [47]), .Z(n3562) );
  CND4X1 U8003 ( .A(n3565), .B(n3564), .C(n3563), .D(n3562), .Z(n1707) );
  CAOR2XL U8004 ( .A(\s1.addr [19]), .B(\s1.dbus_out [60]), .C(n4072), .D(
        \s7.dbus_out [60]), .Z(n3567) );
  CAOR2XL U8005 ( .A(\c1.Breset ), .B(data_stm_d[60]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [60]), .Z(n3566) );
  CANR3X1 U8006 ( .A(n4075), .B(\s6.dbus_out [60]), .C(n3567), .D(n3566), .Z(
        n3576) );
  CND2XL U8007 ( .A(n4098), .B(\s10.dbus_out [60]), .Z(n3571) );
  CANR2XL U8008 ( .A(n4078), .B(\s5.dbus_out [60]), .C(\s4.addr [19]), .D(
        \s4.dbus_out [60]), .Z(n3570) );
  CANR2X1 U8009 ( .A(n4092), .B(\s14.dbus_out [60]), .C(\s12.dbus_out [60]), 
        .D(n4099), .Z(n3569) );
  CND2XL U8010 ( .A(n4101), .B(\s3.dbus_out [60]), .Z(n3568) );
  CAN4X1 U8011 ( .A(n3571), .B(n3570), .C(n3569), .D(n3568), .Z(n3575) );
  CAOR2XL U8012 ( .A(\s9.dbus_out [60]), .B(\s9.addr[7] ), .C(\s0.addr [14]), 
        .D(\s0.dbus_out [60]), .Z(n3572) );
  CANR1XL U8013 ( .A(n4332), .B(\s11.dbus_out [60]), .C(n3572), .Z(n3574) );
  CANR2X1 U8014 ( .A(n4110), .B(\s13.dbus_out [60]), .C(n4085), .D(
        \s8.dbus_out [60]), .Z(n3573) );
  CND4X1 U8015 ( .A(n3576), .B(n3575), .C(n3574), .D(n3573), .Z(n1694) );
  CAOR2X1 U8016 ( .A(n4095), .B(\s1.dbus_out [46]), .C(n4072), .D(
        \s7.dbus_out [46]), .Z(n3578) );
  CAOR2XL U8017 ( .A(\c1.Breset ), .B(data_stm_d[46]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [46]), .Z(n3577) );
  CANR3X1 U8018 ( .A(\s6.addr [17]), .B(\s6.dbus_out [46]), .C(n3578), .D(
        n3577), .Z(n3587) );
  CND2X1 U8019 ( .A(n4098), .B(\s10.dbus_out [46]), .Z(n3582) );
  CANR2X1 U8020 ( .A(n4078), .B(\s5.dbus_out [46]), .C(n4077), .D(
        \s4.dbus_out [46]), .Z(n3581) );
  CANR2X1 U8021 ( .A(n4092), .B(\s14.dbus_out [46]), .C(\s12.dbus_out [46]), 
        .D(n4099), .Z(n3580) );
  CND2XL U8022 ( .A(n4101), .B(\s3.dbus_out [46]), .Z(n3579) );
  CAN4X1 U8023 ( .A(n3582), .B(n3581), .C(n3580), .D(n3579), .Z(n3586) );
  CAOR2XL U8024 ( .A(\s9.dbus_out [46]), .B(n5590), .C(n3940), .D(
        \s0.dbus_out [46]), .Z(n3583) );
  CANR1XL U8025 ( .A(n4108), .B(\s11.dbus_out [46]), .C(n3583), .Z(n3585) );
  CANR2X1 U8026 ( .A(n4110), .B(\s13.dbus_out [46]), .C(n4085), .D(
        \s8.dbus_out [46]), .Z(n3584) );
  CND4X1 U8027 ( .A(n3587), .B(n3586), .C(n3585), .D(n3584), .Z(n1708) );
  CAOR2XL U8028 ( .A(n4090), .B(\s1.dbus_out [57]), .C(n4094), .D(
        \s7.dbus_out [57]), .Z(n3589) );
  CAOR2XL U8029 ( .A(\c1.Breset ), .B(data_stm_d[57]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [57]), .Z(n3588) );
  CANR3X1 U8030 ( .A(\s6.addr [17]), .B(\s6.dbus_out [57]), .C(n3589), .D(
        n3588), .Z(n3598) );
  CND2X1 U8031 ( .A(n4098), .B(\s10.dbus_out [57]), .Z(n3593) );
  CANR2X1 U8032 ( .A(n4078), .B(\s5.dbus_out [57]), .C(n4091), .D(
        \s4.dbus_out [57]), .Z(n3592) );
  CANR2XL U8033 ( .A(n4092), .B(\s14.dbus_out [57]), .C(\s12.dbus_out [57]), 
        .D(n4099), .Z(n3591) );
  CND2XL U8034 ( .A(n4101), .B(\s3.dbus_out [57]), .Z(n3590) );
  CAN4X1 U8035 ( .A(n3593), .B(n3592), .C(n3591), .D(n3590), .Z(n3597) );
  CAOR2XL U8036 ( .A(\s9.dbus_out [57]), .B(\s9.addr [15]), .C(\s0.en ), .D(
        \s0.dbus_out [57]), .Z(n3594) );
  CANR1XL U8037 ( .A(n4108), .B(\s11.dbus_out [57]), .C(n3594), .Z(n3596) );
  CANR2X1 U8038 ( .A(n4110), .B(\s13.dbus_out [57]), .C(n4085), .D(
        \s8.dbus_out [57]), .Z(n3595) );
  CND4X1 U8039 ( .A(n3598), .B(n3597), .C(n3596), .D(n3595), .Z(n1697) );
  CND2XL U8040 ( .A(\s10.en ), .B(\s10.dbus_out [26]), .Z(n3602) );
  CANR2XL U8041 ( .A(n4078), .B(\s5.dbus_out [26]), .C(n4091), .D(
        \s4.dbus_out [26]), .Z(n3601) );
  CANR2XL U8042 ( .A(n4092), .B(\s14.dbus_out [26]), .C(\s12.dbus_out [26]), 
        .D(n4016), .Z(n3600) );
  CND2XL U8043 ( .A(n4101), .B(\s3.dbus_out [26]), .Z(n3599) );
  CAOR2XL U8044 ( .A(\s9.dbus_out [26]), .B(\s9.addr[8] ), .C(\s0.addr [13]), 
        .D(\s0.dbus_out [26]), .Z(n3603) );
  CAOR2X1 U8045 ( .A(n4095), .B(\s1.dbus_out [38]), .C(n4072), .D(
        \s7.dbus_out [38]), .Z(n3605) );
  CAOR2XL U8046 ( .A(\c1.Breset ), .B(data_stm_d[38]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [38]), .Z(n3604) );
  CANR3X1 U8047 ( .A(\s6.addr [17]), .B(\s6.dbus_out [38]), .C(n3605), .D(
        n3604), .Z(n3614) );
  CND2XL U8048 ( .A(\s10.en ), .B(\s10.dbus_out [38]), .Z(n3609) );
  CANR2XL U8049 ( .A(n4078), .B(\s5.dbus_out [38]), .C(n4091), .D(
        \s4.dbus_out [38]), .Z(n3608) );
  CANR2X1 U8050 ( .A(n4092), .B(\s14.dbus_out [38]), .C(\s12.dbus_out [38]), 
        .D(n4099), .Z(n3607) );
  CND2XL U8051 ( .A(n4101), .B(\s3.dbus_out [38]), .Z(n3606) );
  CAN4X1 U8052 ( .A(n3609), .B(n3608), .C(n3607), .D(n3606), .Z(n3613) );
  CAOR2XL U8053 ( .A(\s9.dbus_out [38]), .B(\s9.addr[16] ), .C(n3940), .D(
        \s0.dbus_out [38]), .Z(n3610) );
  CANR1XL U8054 ( .A(n4093), .B(\s11.dbus_out [38]), .C(n3610), .Z(n3612) );
  CANR2X1 U8055 ( .A(n4110), .B(\s13.dbus_out [38]), .C(n4085), .D(
        \s8.dbus_out [38]), .Z(n3611) );
  CND4X1 U8056 ( .A(n3614), .B(n3613), .C(n3612), .D(n3611), .Z(n1716) );
  CAOR2XL U8057 ( .A(n4090), .B(\s1.dbus_out [52]), .C(n4094), .D(
        \s7.dbus_out [52]), .Z(n3616) );
  CAOR2XL U8058 ( .A(\c1.Breset ), .B(data_stm_d[52]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [52]), .Z(n3615) );
  CANR3X1 U8059 ( .A(\s6.addr [17]), .B(\s6.dbus_out [52]), .C(n3616), .D(
        n3615), .Z(n3625) );
  CANR2XL U8060 ( .A(n4078), .B(\s5.dbus_out [52]), .C(n4091), .D(
        \s4.dbus_out [52]), .Z(n3619) );
  CANR2X1 U8061 ( .A(n4092), .B(\s14.dbus_out [52]), .C(\s12.dbus_out [52]), 
        .D(n4099), .Z(n3618) );
  CND2XL U8062 ( .A(n4101), .B(\s3.dbus_out [52]), .Z(n3617) );
  CAN4X1 U8063 ( .A(n3620), .B(n3619), .C(n3618), .D(n3617), .Z(n3624) );
  CAOR2XL U8064 ( .A(\s9.dbus_out [52]), .B(\s9.en ), .C(n4106), .D(
        \s0.dbus_out [52]), .Z(n3621) );
  CANR1XL U8065 ( .A(n4108), .B(\s11.dbus_out [52]), .C(n3621), .Z(n3623) );
  CANR2X1 U8066 ( .A(n4110), .B(\s13.dbus_out [52]), .C(n4109), .D(
        \s8.dbus_out [52]), .Z(n3622) );
  CND4X1 U8067 ( .A(n3625), .B(n3624), .C(n3623), .D(n3622), .Z(n1702) );
  CAOR2XL U8068 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [56]), .C(n4072), .D(
        \s7.dbus_out [56]), .Z(n3627) );
  CAOR2XL U8069 ( .A(\c1.Breset ), .B(data_stm_d[56]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [56]), .Z(n3626) );
  CANR3XL U8070 ( .A(n4062), .B(\s6.dbus_out [56]), .C(n3627), .D(n3626), .Z(
        n3636) );
  CND2XL U8071 ( .A(\s10.en ), .B(\s10.dbus_out [56]), .Z(n3631) );
  CANR2XL U8072 ( .A(n4078), .B(\s5.dbus_out [56]), .C(n4077), .D(
        \s4.dbus_out [56]), .Z(n3630) );
  CANR2XL U8073 ( .A(n4092), .B(\s14.dbus_out [56]), .C(\s12.dbus_out [56]), 
        .D(n4099), .Z(n3629) );
  CND2XL U8074 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [56]), .Z(n3628) );
  CAN4X1 U8075 ( .A(n3631), .B(n3630), .C(n3629), .D(n3628), .Z(n3635) );
  CAOR2XL U8076 ( .A(\s9.dbus_out [56]), .B(\s9.addr[7] ), .C(\s0.en ), .D(
        \s0.dbus_out [56]), .Z(n3632) );
  CANR1XL U8077 ( .A(n4108), .B(\s11.dbus_out [56]), .C(n3632), .Z(n3634) );
  CANR2XL U8078 ( .A(n4110), .B(\s13.dbus_out [56]), .C(n4085), .D(
        \s8.dbus_out [56]), .Z(n3633) );
  CND4X1 U8079 ( .A(n3636), .B(n3635), .C(n3634), .D(n3633), .Z(n1698) );
  CAOR2XL U8080 ( .A(n4090), .B(\s1.dbus_out [37]), .C(n4072), .D(
        \s7.dbus_out [37]), .Z(n3638) );
  CAOR2XL U8081 ( .A(\c1.Breset ), .B(data_stm_d[37]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [37]), .Z(n3637) );
  CANR3X1 U8082 ( .A(n4075), .B(\s6.dbus_out [37]), .C(n3638), .D(n3637), .Z(
        n3647) );
  CND2X1 U8083 ( .A(n4098), .B(\s10.dbus_out [37]), .Z(n3642) );
  CANR2XL U8084 ( .A(n4078), .B(\s5.dbus_out [37]), .C(n4091), .D(
        \s4.dbus_out [37]), .Z(n3641) );
  CANR2XL U8085 ( .A(n4092), .B(\s14.dbus_out [37]), .C(\s12.dbus_out [37]), 
        .D(n1843), .Z(n3640) );
  CND2XL U8086 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [37]), .Z(n3639) );
  CAN4X1 U8087 ( .A(n3642), .B(n3641), .C(n3640), .D(n3639), .Z(n3646) );
  CAOR2XL U8088 ( .A(\s9.dbus_out [37]), .B(\s9.addr[7] ), .C(n4106), .D(
        \s0.dbus_out [37]), .Z(n3643) );
  CANR1XL U8089 ( .A(\s11.dbus_out [37]), .B(n3872), .C(n3643), .Z(n3645) );
  CANR2XL U8090 ( .A(n4110), .B(\s13.dbus_out [37]), .C(\s8.en ), .D(
        \s8.dbus_out [37]), .Z(n3644) );
  CND4X1 U8091 ( .A(n3647), .B(n3646), .C(n3645), .D(n3644), .Z(n1717) );
  CAOR2X1 U8092 ( .A(n4090), .B(\s1.dbus_out [30]), .C(n4094), .D(
        \s7.dbus_out [30]), .Z(n3649) );
  CAOR2XL U8093 ( .A(\c1.Breset ), .B(data_stm_d[30]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [30]), .Z(n3648) );
  CANR3X1 U8094 ( .A(n4075), .B(\s6.dbus_out [30]), .C(n3649), .D(n3648), .Z(
        n3658) );
  CND2X1 U8095 ( .A(n4098), .B(\s10.dbus_out [30]), .Z(n3653) );
  CANR2X1 U8096 ( .A(n4078), .B(\s5.dbus_out [30]), .C(n4077), .D(
        \s4.dbus_out [30]), .Z(n3652) );
  CANR2XL U8097 ( .A(n4100), .B(\s14.dbus_out [30]), .C(\s12.dbus_out [30]), 
        .D(n4099), .Z(n3651) );
  CND2XL U8098 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [30]), .Z(n3650) );
  CAN4X1 U8099 ( .A(n3653), .B(n3652), .C(n3651), .D(n3650), .Z(n3657) );
  CAOR2XL U8100 ( .A(\s9.dbus_out [30]), .B(\s9.addr[8] ), .C(n3963), .D(
        \s0.dbus_out [30]), .Z(n3654) );
  CANR1XL U8101 ( .A(\s11.dbus_out [30]), .B(\s11.addr[17] ), .C(n3654), .Z(
        n3656) );
  CANR2X1 U8102 ( .A(n4110), .B(\s13.dbus_out [30]), .C(n4085), .D(
        \s8.dbus_out [30]), .Z(n3655) );
  CND4X1 U8103 ( .A(n3658), .B(n3657), .C(n3656), .D(n3655), .Z(n1724) );
  CAOR2XL U8104 ( .A(n4090), .B(\s1.dbus_out [44]), .C(n4094), .D(
        \s7.dbus_out [44]), .Z(n3660) );
  CAOR2XL U8105 ( .A(\c1.Breset ), .B(data_stm_d[44]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [44]), .Z(n3659) );
  CANR3X1 U8106 ( .A(n4075), .B(\s6.dbus_out [44]), .C(n3660), .D(n3659), .Z(
        n3669) );
  CND2XL U8107 ( .A(n4098), .B(\s10.dbus_out [44]), .Z(n3664) );
  CANR2XL U8108 ( .A(n4078), .B(\s5.dbus_out [44]), .C(n4091), .D(
        \s4.dbus_out [44]), .Z(n3663) );
  CANR2X1 U8109 ( .A(n4100), .B(\s14.dbus_out [44]), .C(\s12.dbus_out [44]), 
        .D(n4099), .Z(n3662) );
  CND2X1 U8110 ( .A(n4101), .B(\s3.dbus_out [44]), .Z(n3661) );
  CAN4X1 U8111 ( .A(n3664), .B(n3663), .C(n3662), .D(n3661), .Z(n3668) );
  CAOR2XL U8112 ( .A(\s9.dbus_out [44]), .B(n5590), .C(\s0.en ), .D(
        \s0.dbus_out [44]), .Z(n3665) );
  CANR1XL U8113 ( .A(n4108), .B(\s11.dbus_out [44]), .C(n3665), .Z(n3667) );
  CANR2X1 U8114 ( .A(n4110), .B(\s13.dbus_out [44]), .C(n4085), .D(
        \s8.dbus_out [44]), .Z(n3666) );
  CND4X1 U8115 ( .A(n3669), .B(n3668), .C(n3667), .D(n3666), .Z(n1710) );
  CAOR2XL U8116 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [40]), .C(n4072), .D(
        \s7.dbus_out [40]), .Z(n3671) );
  CAOR2XL U8117 ( .A(\c1.Breset ), .B(data_stm_d[40]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [40]), .Z(n3670) );
  CANR3X1 U8118 ( .A(n4075), .B(\s6.dbus_out [40]), .C(n3671), .D(n3670), .Z(
        n3680) );
  CND2X1 U8119 ( .A(n4098), .B(\s10.dbus_out [40]), .Z(n3675) );
  CANR2XL U8120 ( .A(n4078), .B(\s5.dbus_out [40]), .C(n4091), .D(
        \s4.dbus_out [40]), .Z(n3674) );
  CANR2XL U8121 ( .A(n4100), .B(\s14.dbus_out [40]), .C(\s12.dbus_out [40]), 
        .D(n4099), .Z(n3673) );
  CND2X1 U8122 ( .A(n4101), .B(\s3.dbus_out [40]), .Z(n3672) );
  CAN4X1 U8123 ( .A(n3675), .B(n3674), .C(n3673), .D(n3672), .Z(n3679) );
  CAOR2XL U8124 ( .A(\s9.dbus_out [40]), .B(\s9.addr[8] ), .C(n4083), .D(
        \s0.dbus_out [40]), .Z(n3676) );
  CANR1XL U8125 ( .A(n4108), .B(\s11.dbus_out [40]), .C(n3676), .Z(n3678) );
  CANR2XL U8126 ( .A(n4110), .B(\s13.dbus_out [40]), .C(n4109), .D(
        \s8.dbus_out [40]), .Z(n3677) );
  CND4X1 U8127 ( .A(n3680), .B(n3679), .C(n3678), .D(n3677), .Z(n1714) );
  CAOR2X1 U8128 ( .A(n4090), .B(\s1.dbus_out [3]), .C(n4094), .D(
        \s7.dbus_out [3]), .Z(n3682) );
  CAOR2XL U8129 ( .A(\c1.Breset ), .B(data_stm_d[3]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [3]), .Z(n3681) );
  CANR3X1 U8130 ( .A(\s6.addr [17]), .B(\s6.dbus_out [3]), .C(n3682), .D(n3681), .Z(n3691) );
  CND2XL U8131 ( .A(n4050), .B(\s10.dbus_out [3]), .Z(n3686) );
  CANR2XL U8132 ( .A(n4078), .B(\s5.dbus_out [3]), .C(n4091), .D(
        \s4.dbus_out [3]), .Z(n3685) );
  CANR2X1 U8133 ( .A(n4100), .B(\s14.dbus_out [3]), .C(\s12.dbus_out [3]), .D(
        n4099), .Z(n3684) );
  CND2X1 U8134 ( .A(n4101), .B(\s3.dbus_out [3]), .Z(n3683) );
  CAN4X1 U8135 ( .A(n3686), .B(n3685), .C(n3684), .D(n3683), .Z(n3690) );
  CAOR2XL U8136 ( .A(\s9.dbus_out [3]), .B(\s9.addr[7] ), .C(n3940), .D(
        \s0.dbus_out [3]), .Z(n3687) );
  CANR1XL U8137 ( .A(n4093), .B(\s11.dbus_out [3]), .C(n3687), .Z(n3689) );
  CANR2XL U8138 ( .A(n4110), .B(\s13.dbus_out [3]), .C(\s8.addr[15] ), .D(
        \s8.dbus_out [3]), .Z(n3688) );
  CND4X1 U8139 ( .A(n3691), .B(n3690), .C(n3689), .D(n3688), .Z(n1751) );
  CAOR2X1 U8140 ( .A(n4090), .B(\s1.dbus_out [12]), .C(n4072), .D(
        \s7.dbus_out [12]), .Z(n3693) );
  CAOR2XL U8141 ( .A(\c1.Breset ), .B(data_stm_d[12]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [12]), .Z(n3692) );
  CANR3X1 U8142 ( .A(\s6.addr [17]), .B(\s6.dbus_out [12]), .C(n3693), .D(
        n3692), .Z(n3702) );
  CND2X1 U8143 ( .A(n4098), .B(\s10.dbus_out [12]), .Z(n3697) );
  CANR2XL U8144 ( .A(n4078), .B(\s5.dbus_out [12]), .C(n4091), .D(
        \s4.dbus_out [12]), .Z(n3696) );
  CANR2XL U8145 ( .A(n4092), .B(\s14.dbus_out [12]), .C(\s12.dbus_out [12]), 
        .D(n1840), .Z(n3695) );
  CND2XL U8146 ( .A(\s3.addr [18]), .B(\s3.dbus_out [12]), .Z(n3694) );
  CAN4X1 U8147 ( .A(n3697), .B(n3696), .C(n3695), .D(n3694), .Z(n3701) );
  CAOR2XL U8148 ( .A(\s9.dbus_out [12]), .B(\s9.addr[16] ), .C(\s0.addr [13]), 
        .D(\s0.dbus_out [12]), .Z(n3698) );
  CANR1XL U8149 ( .A(n4093), .B(\s11.dbus_out [12]), .C(n3698), .Z(n3700) );
  CANR2XL U8150 ( .A(n4110), .B(\s13.dbus_out [12]), .C(\s8.dbus_out [12]), 
        .D(n4109), .Z(n3699) );
  CND4X1 U8151 ( .A(n3702), .B(n3701), .C(n3700), .D(n3699), .Z(n1742) );
  CAOR2X1 U8152 ( .A(n4090), .B(\s1.dbus_out [13]), .C(n4072), .D(
        \s7.dbus_out [13]), .Z(n3704) );
  CAOR2XL U8153 ( .A(\c1.Breset ), .B(data_stm_d[13]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [13]), .Z(n3703) );
  CANR3X1 U8154 ( .A(\s6.addr [17]), .B(\s6.dbus_out [13]), .C(n3704), .D(
        n3703), .Z(n3714) );
  CNR2IX1 U8155 ( .B(\s10.dbus_out [13]), .A(n4076), .Z(n3705) );
  CIVX2 U8156 ( .A(n3705), .Z(n3709) );
  CANR2XL U8157 ( .A(n4078), .B(\s5.dbus_out [13]), .C(n4091), .D(
        \s4.dbus_out [13]), .Z(n3708) );
  CANR2X1 U8158 ( .A(n4100), .B(\s14.dbus_out [13]), .C(\s12.dbus_out [13]), 
        .D(n4099), .Z(n3707) );
  CND2XL U8159 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [13]), .Z(n3706) );
  CAN4X1 U8160 ( .A(n3709), .B(n3708), .C(n3707), .D(n3706), .Z(n3713) );
  CAOR2XL U8161 ( .A(\s9.dbus_out [13]), .B(\s9.addr[8] ), .C(n4106), .D(
        \s0.dbus_out [13]), .Z(n3710) );
  CANR1XL U8162 ( .A(n4093), .B(\s11.dbus_out [13]), .C(n3710), .Z(n3712) );
  CANR2X1 U8163 ( .A(n4110), .B(\s13.dbus_out [13]), .C(n4085), .D(
        \s8.dbus_out [13]), .Z(n3711) );
  CND4X1 U8164 ( .A(n3714), .B(n3713), .C(n3712), .D(n3711), .Z(n1741) );
  CAOR2XL U8165 ( .A(n4090), .B(\s1.dbus_out [2]), .C(n4094), .D(
        \s7.dbus_out [2]), .Z(n3716) );
  CAOR2XL U8166 ( .A(\c1.Breset ), .B(data_stm_d[2]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [2]), .Z(n3715) );
  CANR3XL U8167 ( .A(\s6.en ), .B(\s6.dbus_out [2]), .C(n3716), .D(n3715), .Z(
        n3725) );
  CND2X1 U8168 ( .A(n4098), .B(\s10.dbus_out [2]), .Z(n3720) );
  CANR2XL U8169 ( .A(n4078), .B(\s5.dbus_out [2]), .C(n4091), .D(
        \s4.dbus_out [2]), .Z(n3719) );
  CANR2XL U8170 ( .A(n4100), .B(\s14.dbus_out [2]), .C(\s12.dbus_out [2]), .D(
        n4099), .Z(n3718) );
  CND2X1 U8171 ( .A(n4101), .B(\s3.dbus_out [2]), .Z(n3717) );
  CAN4X1 U8172 ( .A(n3720), .B(n3719), .C(n3718), .D(n3717), .Z(n3724) );
  CAOR2XL U8173 ( .A(\s9.dbus_out [2]), .B(n5590), .C(n4106), .D(
        \s0.dbus_out [2]), .Z(n3721) );
  CANR1XL U8174 ( .A(n4108), .B(\s11.dbus_out [2]), .C(n3721), .Z(n3723) );
  CANR2X1 U8175 ( .A(n4110), .B(\s13.dbus_out [2]), .C(n4085), .D(
        \s8.dbus_out [2]), .Z(n3722) );
  CND4X1 U8176 ( .A(n3725), .B(n3724), .C(n3723), .D(n3722), .Z(n1752) );
  CAOR2XL U8177 ( .A(n4090), .B(\s1.dbus_out [7]), .C(n4094), .D(
        \s7.dbus_out [7]), .Z(n3727) );
  CAOR2XL U8178 ( .A(\c1.Breset ), .B(data_stm_d[7]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [7]), .Z(n3726) );
  CANR3X1 U8179 ( .A(\s6.addr [17]), .B(\s6.dbus_out [7]), .C(n3727), .D(n3726), .Z(n3736) );
  CND2XL U8180 ( .A(\s10.addr[9] ), .B(\s10.dbus_out [7]), .Z(n3731) );
  CANR2XL U8181 ( .A(n4078), .B(\s5.dbus_out [7]), .C(n4091), .D(
        \s4.dbus_out [7]), .Z(n3730) );
  CANR2XL U8182 ( .A(n4092), .B(\s14.dbus_out [7]), .C(\s12.dbus_out [7]), .D(
        n4099), .Z(n3729) );
  CND2X1 U8183 ( .A(n4101), .B(\s3.dbus_out [7]), .Z(n3728) );
  CAN4X1 U8184 ( .A(n3731), .B(n3730), .C(n3729), .D(n3728), .Z(n3735) );
  CAOR2XL U8185 ( .A(\s9.dbus_out [7]), .B(\s9.addr[7] ), .C(n3963), .D(
        \s0.dbus_out [7]), .Z(n3732) );
  CANR1XL U8186 ( .A(n4108), .B(\s11.dbus_out [7]), .C(n3732), .Z(n3734) );
  CANR2X1 U8187 ( .A(n4110), .B(\s13.dbus_out [7]), .C(n4085), .D(
        \s8.dbus_out [7]), .Z(n3733) );
  CND4X1 U8188 ( .A(n3736), .B(n3735), .C(n3734), .D(n3733), .Z(n1747) );
  CAOR2XL U8189 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [5]), .C(n4094), .D(
        \s7.dbus_out [5]), .Z(n3738) );
  CAOR2XL U8190 ( .A(\c1.Breset ), .B(data_stm_d[5]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [5]), .Z(n3737) );
  CANR3XL U8191 ( .A(n4062), .B(\s6.dbus_out [5]), .C(n3738), .D(n3737), .Z(
        n3747) );
  CND2XL U8192 ( .A(n4050), .B(\s10.dbus_out [5]), .Z(n3742) );
  CANR2XL U8193 ( .A(n4078), .B(\s5.dbus_out [5]), .C(n4091), .D(
        \s4.dbus_out [5]), .Z(n3741) );
  CANR2X1 U8194 ( .A(n4100), .B(\s14.dbus_out [5]), .C(\s12.dbus_out [5]), .D(
        n4099), .Z(n3740) );
  CND2X1 U8195 ( .A(n4101), .B(\s3.dbus_out [5]), .Z(n3739) );
  CAN4X1 U8196 ( .A(n3742), .B(n3741), .C(n3740), .D(n3739), .Z(n3746) );
  CAOR2XL U8197 ( .A(\s9.dbus_out [5]), .B(\s9.addr[16] ), .C(n3963), .D(
        \s0.dbus_out [5]), .Z(n3743) );
  CANR1XL U8198 ( .A(n4093), .B(\s11.dbus_out [5]), .C(n3743), .Z(n3745) );
  CANR2XL U8199 ( .A(n4110), .B(\s13.dbus_out [5]), .C(\s8.en ), .D(
        \s8.dbus_out [5]), .Z(n3744) );
  CND4X1 U8200 ( .A(n3747), .B(n3746), .C(n3745), .D(n3744), .Z(n1749) );
  CND2XL U8201 ( .A(\s10.en ), .B(\s10.dbus_out [11]), .Z(n3751) );
  CANR2XL U8202 ( .A(n4078), .B(\s5.dbus_out [11]), .C(n4091), .D(
        \s4.dbus_out [11]), .Z(n3750) );
  CANR2XL U8203 ( .A(n4092), .B(\s14.dbus_out [11]), .C(\s12.dbus_out [11]), 
        .D(n1840), .Z(n3749) );
  CND2XL U8204 ( .A(n4101), .B(\s3.dbus_out [11]), .Z(n3748) );
  CAN4X1 U8205 ( .A(n3751), .B(n3750), .C(n3749), .D(n3748), .Z(n3755) );
  CAOR2XL U8206 ( .A(\s9.dbus_out [11]), .B(\s9.addr[8] ), .C(n3975), .D(
        \s0.dbus_out [11]), .Z(n3752) );
  CANR1XL U8207 ( .A(n4093), .B(\s11.dbus_out [11]), .C(n3752), .Z(n3754) );
  CANR2XL U8208 ( .A(n4110), .B(\s13.dbus_out [11]), .C(n4085), .D(
        \s8.dbus_out [11]), .Z(n3753) );
  CND4X1 U8209 ( .A(n3756), .B(n3755), .C(n3754), .D(n3753), .Z(n1743) );
  CAOR2X1 U8210 ( .A(n4090), .B(\s1.dbus_out [6]), .C(n4094), .D(
        \s7.dbus_out [6]), .Z(n3758) );
  CAOR2XL U8211 ( .A(\c1.Breset ), .B(data_stm_d[6]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [6]), .Z(n3757) );
  CANR3X1 U8212 ( .A(\s6.addr [17]), .B(\s6.dbus_out [6]), .C(n3758), .D(n3757), .Z(n3767) );
  CND2X1 U8213 ( .A(n4098), .B(\s10.dbus_out [6]), .Z(n3762) );
  CANR2XL U8214 ( .A(n4078), .B(\s5.dbus_out [6]), .C(\s4.addr [19]), .D(
        \s4.dbus_out [6]), .Z(n3761) );
  CANR2X1 U8215 ( .A(n4100), .B(\s14.dbus_out [6]), .C(\s12.dbus_out [6]), .D(
        n4099), .Z(n3760) );
  CND2XL U8216 ( .A(\s3.addr [18]), .B(\s3.dbus_out [6]), .Z(n3759) );
  CAN4X1 U8217 ( .A(n3762), .B(n3761), .C(n3760), .D(n3759), .Z(n3766) );
  CAOR2XL U8218 ( .A(\s9.dbus_out [6]), .B(\s9.en ), .C(\s0.addr [12]), .D(
        \s0.dbus_out [6]), .Z(n3763) );
  CANR1XL U8219 ( .A(n4093), .B(\s11.dbus_out [6]), .C(n3763), .Z(n3765) );
  CANR2XL U8220 ( .A(n4110), .B(\s13.dbus_out [6]), .C(\s8.en ), .D(
        \s8.dbus_out [6]), .Z(n3764) );
  CND4X1 U8221 ( .A(n3767), .B(n3766), .C(n3765), .D(n3764), .Z(n1748) );
  CND2XL U8222 ( .A(\s10.en ), .B(\s10.dbus_out [9]), .Z(n3771) );
  CANR2XL U8223 ( .A(n4078), .B(\s5.dbus_out [9]), .C(n4091), .D(
        \s4.dbus_out [9]), .Z(n3770) );
  CANR2XL U8224 ( .A(\s14.addr[16] ), .B(\s14.dbus_out [9]), .C(
        \s12.dbus_out [9]), .D(n1840), .Z(n3769) );
  CND2XL U8225 ( .A(n4101), .B(\s3.dbus_out [9]), .Z(n3768) );
  CAN4X1 U8226 ( .A(n3771), .B(n3770), .C(n3769), .D(n3768), .Z(n3775) );
  CAOR2XL U8227 ( .A(\s9.dbus_out [9]), .B(\s9.addr[8] ), .C(n3963), .D(
        \s0.dbus_out [9]), .Z(n3772) );
  CANR1XL U8228 ( .A(n4108), .B(\s11.dbus_out [9]), .C(n3772), .Z(n3774) );
  CANR2X1 U8229 ( .A(n4110), .B(\s13.dbus_out [9]), .C(n4109), .D(
        \s8.dbus_out [9]), .Z(n3773) );
  CND4X1 U8230 ( .A(n3776), .B(n3775), .C(n3774), .D(n3773), .Z(n1745) );
  CAOR2XL U8231 ( .A(\s1.addr [19]), .B(\s1.dbus_out [10]), .C(n4094), .D(
        \s7.dbus_out [10]), .Z(n3778) );
  CAOR2XL U8232 ( .A(\c1.Breset ), .B(data_stm_d[10]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [10]), .Z(n3777) );
  CANR3X1 U8233 ( .A(\s6.addr [17]), .B(\s6.dbus_out [10]), .C(n3778), .D(
        n3777), .Z(n3787) );
  CND2XL U8234 ( .A(\s10.addr[9] ), .B(\s10.dbus_out [10]), .Z(n3782) );
  CANR2XL U8235 ( .A(n4078), .B(\s5.dbus_out [10]), .C(n4077), .D(
        \s4.dbus_out [10]), .Z(n3781) );
  CANR2X1 U8236 ( .A(n4092), .B(\s14.dbus_out [10]), .C(\s12.dbus_out [10]), 
        .D(n4099), .Z(n3780) );
  CND2XL U8237 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [10]), .Z(n3779) );
  CAN4X1 U8238 ( .A(n3782), .B(n3781), .C(n3780), .D(n3779), .Z(n3786) );
  CAOR2XL U8239 ( .A(\s9.dbus_out [10]), .B(\s9.addr[16] ), .C(\s0.addr [14]), 
        .D(\s0.dbus_out [10]), .Z(n3783) );
  CANR1XL U8240 ( .A(\s11.en ), .B(\s11.dbus_out [10]), .C(n3783), .Z(n3785)
         );
  CANR2XL U8241 ( .A(n4110), .B(\s13.dbus_out [10]), .C(\s8.addr[15] ), .D(
        \s8.dbus_out [10]), .Z(n3784) );
  CND4X1 U8242 ( .A(n3787), .B(n3786), .C(n3785), .D(n3784), .Z(n1744) );
  CAOR2XL U8243 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [4]), .C(n4072), .D(
        \s7.dbus_out [4]), .Z(n3789) );
  CAOR2XL U8244 ( .A(\c1.Breset ), .B(data_stm_d[4]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [4]), .Z(n3788) );
  CANR3X1 U8245 ( .A(\s6.addr [17]), .B(\s6.dbus_out [4]), .C(n3789), .D(n3788), .Z(n3798) );
  CND2X1 U8246 ( .A(n4098), .B(\s10.dbus_out [4]), .Z(n3793) );
  CANR2X1 U8247 ( .A(n4078), .B(\s5.dbus_out [4]), .C(n4077), .D(
        \s4.dbus_out [4]), .Z(n3792) );
  CANR2XL U8248 ( .A(\s14.addr [11]), .B(\s14.dbus_out [4]), .C(
        \s12.dbus_out [4]), .D(n4099), .Z(n3791) );
  CND2X1 U8249 ( .A(n4101), .B(\s3.dbus_out [4]), .Z(n3790) );
  CAN4X1 U8250 ( .A(n3793), .B(n3792), .C(n3791), .D(n3790), .Z(n3797) );
  CAOR2XL U8251 ( .A(\s9.dbus_out [4]), .B(\s9.addr[7] ), .C(n3975), .D(
        \s0.dbus_out [4]), .Z(n3794) );
  CANR1XL U8252 ( .A(n4108), .B(\s11.dbus_out [4]), .C(n3794), .Z(n3796) );
  CANR2XL U8253 ( .A(n4110), .B(\s13.dbus_out [4]), .C(\s8.dbus_out [4]), .D(
        n4085), .Z(n3795) );
  CND4X1 U8254 ( .A(n3798), .B(n3797), .C(n3796), .D(n3795), .Z(n1750) );
  CAOR2XL U8255 ( .A(\s1.addr [19]), .B(\s1.dbus_out [51]), .C(n4072), .D(
        \s7.dbus_out [51]), .Z(n3800) );
  CAOR2XL U8256 ( .A(\c1.Breset ), .B(data_stm_d[51]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [51]), .Z(n3799) );
  CANR3X1 U8257 ( .A(\s6.addr [17]), .B(\s6.dbus_out [51]), .C(n3800), .D(
        n3799), .Z(n3809) );
  CND2XL U8258 ( .A(n4098), .B(\s10.dbus_out [51]), .Z(n3804) );
  CANR2XL U8259 ( .A(n4078), .B(\s5.dbus_out [51]), .C(\s4.addr [19]), .D(
        \s4.dbus_out [51]), .Z(n3803) );
  CANR2XL U8260 ( .A(n4100), .B(\s14.dbus_out [51]), .C(\s12.dbus_out [51]), 
        .D(n1843), .Z(n3802) );
  CND2XL U8261 ( .A(n4101), .B(\s3.dbus_out [51]), .Z(n3801) );
  CAN4X1 U8262 ( .A(n3804), .B(n3803), .C(n3802), .D(n3801), .Z(n3808) );
  CAOR2XL U8263 ( .A(\s9.dbus_out [51]), .B(\s9.addr[8] ), .C(n3963), .D(
        \s0.dbus_out [51]), .Z(n3805) );
  CANR1XL U8264 ( .A(\s11.en ), .B(\s11.dbus_out [51]), .C(n3805), .Z(n3807)
         );
  CANR2XL U8265 ( .A(n4110), .B(\s13.dbus_out [51]), .C(\s8.en ), .D(
        \s8.dbus_out [51]), .Z(n3806) );
  CND4X1 U8266 ( .A(n3809), .B(n3808), .C(n3807), .D(n3806), .Z(n1703) );
  CAOR2XL U8267 ( .A(\s1.addr [19]), .B(\s1.dbus_out [45]), .C(\s7.addr[16] ), 
        .D(\s7.dbus_out [45]), .Z(n3811) );
  CAOR2XL U8268 ( .A(\c1.Breset ), .B(data_stm_d[45]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [45]), .Z(n3810) );
  CANR3X1 U8269 ( .A(n4075), .B(\s6.dbus_out [45]), .C(n3811), .D(n3810), .Z(
        n3820) );
  CND2XL U8270 ( .A(n4098), .B(\s10.dbus_out [45]), .Z(n3815) );
  CANR2X1 U8271 ( .A(n4078), .B(\s5.dbus_out [45]), .C(n4091), .D(
        \s4.dbus_out [45]), .Z(n3814) );
  CANR2X1 U8272 ( .A(n4092), .B(\s14.dbus_out [45]), .C(\s12.dbus_out [45]), 
        .D(n4099), .Z(n3813) );
  CND2X1 U8273 ( .A(n4101), .B(\s3.dbus_out [45]), .Z(n3812) );
  CAN4X1 U8274 ( .A(n3815), .B(n3814), .C(n3813), .D(n3812), .Z(n3819) );
  CAOR2XL U8275 ( .A(\s9.dbus_out [45]), .B(\s9.addr[16] ), .C(\s0.addr [12]), 
        .D(\s0.dbus_out [45]), .Z(n3816) );
  CANR1XL U8276 ( .A(n4108), .B(\s11.dbus_out [45]), .C(n3816), .Z(n3818) );
  CANR2XL U8277 ( .A(n4110), .B(\s13.dbus_out [45]), .C(\s8.en ), .D(
        \s8.dbus_out [45]), .Z(n3817) );
  CND4X1 U8278 ( .A(n3820), .B(n3819), .C(n3818), .D(n3817), .Z(n1709) );
  CAOR2X1 U8279 ( .A(n4090), .B(\s1.dbus_out [55]), .C(n4072), .D(
        \s7.dbus_out [55]), .Z(n3822) );
  CAOR2XL U8280 ( .A(\c1.Breset ), .B(data_stm_d[55]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [55]), .Z(n3821) );
  CANR3X1 U8281 ( .A(\s6.addr [17]), .B(\s6.dbus_out [55]), .C(n3822), .D(
        n3821), .Z(n3831) );
  CND2XL U8282 ( .A(n4098), .B(\s10.dbus_out [55]), .Z(n3826) );
  CANR2XL U8283 ( .A(n4078), .B(\s5.dbus_out [55]), .C(n4077), .D(
        \s4.dbus_out [55]), .Z(n3825) );
  CANR2XL U8284 ( .A(n4092), .B(\s14.dbus_out [55]), .C(\s12.dbus_out [55]), 
        .D(n1843), .Z(n3824) );
  CND2XL U8285 ( .A(n4101), .B(\s3.dbus_out [55]), .Z(n3823) );
  CAN4X1 U8286 ( .A(n3826), .B(n3825), .C(n3824), .D(n3823), .Z(n3830) );
  CAOR2XL U8287 ( .A(\s9.dbus_out [55]), .B(\s9.addr[8] ), .C(n4106), .D(
        \s0.dbus_out [55]), .Z(n3827) );
  CANR1XL U8288 ( .A(n4093), .B(\s11.dbus_out [55]), .C(n3827), .Z(n3829) );
  CANR2XL U8289 ( .A(n4110), .B(\s13.dbus_out [55]), .C(\s8.en ), .D(
        \s8.dbus_out [55]), .Z(n3828) );
  CND4X1 U8290 ( .A(n3831), .B(n3830), .C(n3829), .D(n3828), .Z(n1699) );
  CAOR2X1 U8291 ( .A(n4090), .B(\s1.dbus_out [49]), .C(n4094), .D(
        \s7.dbus_out [49]), .Z(n3833) );
  CAOR2XL U8292 ( .A(\c1.Breset ), .B(data_stm_d[49]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [49]), .Z(n3832) );
  CANR3X1 U8293 ( .A(\s6.addr [17]), .B(\s6.dbus_out [49]), .C(n3833), .D(
        n3832), .Z(n3842) );
  CND2X1 U8294 ( .A(n4098), .B(\s10.dbus_out [49]), .Z(n3837) );
  CANR2XL U8295 ( .A(n4078), .B(\s5.dbus_out [49]), .C(n4077), .D(
        \s4.dbus_out [49]), .Z(n3836) );
  CANR2XL U8296 ( .A(n4100), .B(\s14.dbus_out [49]), .C(\s12.dbus_out [49]), 
        .D(n1843), .Z(n3835) );
  CND2XL U8297 ( .A(n4101), .B(\s3.dbus_out [49]), .Z(n3834) );
  CAN4X1 U8298 ( .A(n3837), .B(n3836), .C(n3835), .D(n3834), .Z(n3841) );
  CAOR2XL U8299 ( .A(\s9.dbus_out [49]), .B(\s9.addr[16] ), .C(n3975), .D(
        \s0.dbus_out [49]), .Z(n3838) );
  CANR1XL U8300 ( .A(n4108), .B(\s11.dbus_out [49]), .C(n3838), .Z(n3840) );
  CANR2X1 U8301 ( .A(n4110), .B(\s13.dbus_out [49]), .C(n4085), .D(
        \s8.dbus_out [49]), .Z(n3839) );
  CND4X1 U8302 ( .A(n3842), .B(n3841), .C(n3840), .D(n3839), .Z(n1705) );
  CAOR2XL U8303 ( .A(n4090), .B(\s1.dbus_out [16]), .C(n4094), .D(
        \s7.dbus_out [16]), .Z(n3844) );
  CAOR2XL U8304 ( .A(\c1.Breset ), .B(data_stm_d[16]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [16]), .Z(n3843) );
  CANR3X1 U8305 ( .A(n4075), .B(\s6.dbus_out [16]), .C(n3844), .D(n3843), .Z(
        n3853) );
  CND2XL U8306 ( .A(n4050), .B(\s10.dbus_out [16]), .Z(n3848) );
  CANR2XL U8307 ( .A(n4078), .B(\s5.dbus_out [16]), .C(n4077), .D(
        \s4.dbus_out [16]), .Z(n3847) );
  CANR2X1 U8308 ( .A(n4100), .B(\s14.dbus_out [16]), .C(\s12.dbus_out [16]), 
        .D(n4099), .Z(n3846) );
  CND2XL U8309 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [16]), .Z(n3845) );
  CAN4X1 U8310 ( .A(n3848), .B(n3847), .C(n3846), .D(n3845), .Z(n3852) );
  CAOR2XL U8311 ( .A(\s9.dbus_out [16]), .B(\s9.addr [15]), .C(n3940), .D(
        \s0.dbus_out [16]), .Z(n3849) );
  CANR1XL U8312 ( .A(\s11.en ), .B(\s11.dbus_out [16]), .C(n3849), .Z(n3851)
         );
  CANR2XL U8313 ( .A(n4110), .B(\s13.dbus_out [16]), .C(n4085), .D(
        \s8.dbus_out [16]), .Z(n3850) );
  CND4X1 U8314 ( .A(n3853), .B(n3852), .C(n3851), .D(n3850), .Z(n1738) );
  CAOR2X1 U8315 ( .A(n4090), .B(\s1.dbus_out [63]), .C(n4094), .D(
        \s7.dbus_out [63]), .Z(n3855) );
  CAOR2XL U8316 ( .A(\c1.Breset ), .B(data_stm_d[63]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [63]), .Z(n3854) );
  CANR3X1 U8317 ( .A(n4075), .B(\s6.dbus_out [63]), .C(n3855), .D(n3854), .Z(
        n3864) );
  CND2XL U8318 ( .A(n4050), .B(\s10.dbus_out [63]), .Z(n3859) );
  CANR2XL U8319 ( .A(n4078), .B(\s5.dbus_out [63]), .C(n4091), .D(
        \s4.dbus_out [63]), .Z(n3858) );
  CANR2XL U8320 ( .A(n4100), .B(\s14.dbus_out [63]), .C(\s12.dbus_out [63]), 
        .D(n4099), .Z(n3857) );
  CND2XL U8321 ( .A(\s3.addr [18]), .B(\s3.dbus_out [63]), .Z(n3856) );
  CAN4X1 U8322 ( .A(n3859), .B(n3858), .C(n3857), .D(n3856), .Z(n3863) );
  CAOR2XL U8323 ( .A(\s9.dbus_out [63]), .B(\s9.addr[8] ), .C(n3975), .D(
        \s0.dbus_out [63]), .Z(n3860) );
  CANR1XL U8324 ( .A(n4093), .B(\s11.dbus_out [63]), .C(n3860), .Z(n3862) );
  CANR2XL U8325 ( .A(n4110), .B(\s13.dbus_out [63]), .C(n4109), .D(
        \s8.dbus_out [63]), .Z(n3861) );
  CND4X1 U8326 ( .A(n3864), .B(n3863), .C(n3862), .D(n3861), .Z(n1691) );
  CAOR2X1 U8327 ( .A(n4090), .B(\s1.dbus_out [50]), .C(n4072), .D(
        \s7.dbus_out [50]), .Z(n3866) );
  CAOR2XL U8328 ( .A(\c1.Breset ), .B(data_stm_d[50]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [50]), .Z(n3865) );
  CANR3X1 U8329 ( .A(n4075), .B(\s6.dbus_out [50]), .C(n3866), .D(n3865), .Z(
        n3876) );
  CND2XL U8330 ( .A(n4050), .B(\s10.dbus_out [50]), .Z(n3870) );
  CANR2XL U8331 ( .A(n4078), .B(\s5.dbus_out [50]), .C(\s4.addr [19]), .D(
        \s4.dbus_out [50]), .Z(n3869) );
  CANR2X1 U8332 ( .A(n4100), .B(\s14.dbus_out [50]), .C(\s12.dbus_out [50]), 
        .D(n4099), .Z(n3868) );
  CND2XL U8333 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [50]), .Z(n3867) );
  CAN4X1 U8334 ( .A(n3870), .B(n3869), .C(n3868), .D(n3867), .Z(n3875) );
  CAOR2XL U8335 ( .A(\s9.dbus_out [50]), .B(\s9.addr[7] ), .C(n3975), .D(
        \s0.dbus_out [50]), .Z(n3871) );
  CANR1XL U8336 ( .A(\s11.dbus_out [50]), .B(n3872), .C(n3871), .Z(n3874) );
  CANR2X1 U8337 ( .A(n4110), .B(\s13.dbus_out [50]), .C(n4085), .D(
        \s8.dbus_out [50]), .Z(n3873) );
  CND4X1 U8338 ( .A(n3876), .B(n3875), .C(n3874), .D(n3873), .Z(n1704) );
  CAOR2XL U8339 ( .A(\s1.addr [19]), .B(\s1.dbus_out [54]), .C(n4094), .D(
        \s7.dbus_out [54]), .Z(n3878) );
  CAOR2XL U8340 ( .A(\c1.Breset ), .B(data_stm_d[54]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [54]), .Z(n3877) );
  CANR3X1 U8341 ( .A(n4075), .B(\s6.dbus_out [54]), .C(n3878), .D(n3877), .Z(
        n3887) );
  CANR2XL U8342 ( .A(n4078), .B(\s5.dbus_out [54]), .C(n4077), .D(
        \s4.dbus_out [54]), .Z(n3881) );
  CANR2XL U8343 ( .A(n4092), .B(\s14.dbus_out [54]), .C(\s12.dbus_out [54]), 
        .D(n1843), .Z(n3880) );
  CND2XL U8344 ( .A(n4101), .B(\s3.dbus_out [54]), .Z(n3879) );
  CAN4X1 U8345 ( .A(n3882), .B(n3881), .C(n3880), .D(n3879), .Z(n3886) );
  CAOR2XL U8346 ( .A(\s9.dbus_out [54]), .B(n5590), .C(n3963), .D(
        \s0.dbus_out [54]), .Z(n3883) );
  CANR1XL U8347 ( .A(n4108), .B(\s11.dbus_out [54]), .C(n3883), .Z(n3885) );
  CANR2X1 U8348 ( .A(n4110), .B(\s13.dbus_out [54]), .C(n4085), .D(
        \s8.dbus_out [54]), .Z(n3884) );
  CND4X1 U8349 ( .A(n3887), .B(n3886), .C(n3885), .D(n3884), .Z(n1700) );
  CAOR2X1 U8350 ( .A(n4095), .B(\s1.dbus_out [31]), .C(n4072), .D(
        \s7.dbus_out [31]), .Z(n3889) );
  CAOR2XL U8351 ( .A(\c1.Breset ), .B(data_stm_d[31]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [31]), .Z(n3888) );
  CANR3XL U8352 ( .A(n4062), .B(\s6.dbus_out [31]), .C(n3889), .D(n3888), .Z(
        n3898) );
  CND2X1 U8353 ( .A(n4098), .B(\s10.dbus_out [31]), .Z(n3893) );
  CANR2XL U8354 ( .A(n4078), .B(\s5.dbus_out [31]), .C(n4077), .D(
        \s4.dbus_out [31]), .Z(n3892) );
  CANR2X1 U8355 ( .A(n4092), .B(\s14.dbus_out [31]), .C(\s12.dbus_out [31]), 
        .D(n4099), .Z(n3891) );
  CND2XL U8356 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [31]), .Z(n3890) );
  CAN4X1 U8357 ( .A(n3893), .B(n3892), .C(n3891), .D(n3890), .Z(n3897) );
  CAOR2XL U8358 ( .A(\s9.dbus_out [31]), .B(\s9.addr [15]), .C(n4083), .D(
        \s0.dbus_out [31]), .Z(n3894) );
  CANR1XL U8359 ( .A(n4108), .B(\s11.dbus_out [31]), .C(n3894), .Z(n3896) );
  CANR2X1 U8360 ( .A(n4110), .B(\s13.dbus_out [31]), .C(n4085), .D(
        \s8.dbus_out [31]), .Z(n3895) );
  CND4X1 U8361 ( .A(n3898), .B(n3897), .C(n3896), .D(n3895), .Z(n1723) );
  CAOR2XL U8362 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [53]), .C(n4094), .D(
        \s7.dbus_out [53]), .Z(n3900) );
  CAOR2XL U8363 ( .A(\c1.Breset ), .B(data_stm_d[53]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [53]), .Z(n3899) );
  CANR3X1 U8364 ( .A(n4075), .B(\s6.dbus_out [53]), .C(n3900), .D(n3899), .Z(
        n3910) );
  CNR2IX1 U8365 ( .B(\s10.dbus_out [53]), .A(n4076), .Z(n3901) );
  CIVX2 U8366 ( .A(n3901), .Z(n3905) );
  CANR2XL U8367 ( .A(n4078), .B(\s5.dbus_out [53]), .C(\s4.addr [19]), .D(
        \s4.dbus_out [53]), .Z(n3904) );
  CANR2X1 U8368 ( .A(n4092), .B(\s14.dbus_out [53]), .C(\s12.dbus_out [53]), 
        .D(n4099), .Z(n3903) );
  CND2XL U8369 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [53]), .Z(n3902) );
  CAN4X1 U8370 ( .A(n3905), .B(n3904), .C(n3903), .D(n3902), .Z(n3909) );
  CAOR2XL U8371 ( .A(\s9.dbus_out [53]), .B(\s9.addr[16] ), .C(n4106), .D(
        \s0.dbus_out [53]), .Z(n3906) );
  CANR1XL U8372 ( .A(n4108), .B(\s11.dbus_out [53]), .C(n3906), .Z(n3908) );
  CANR2X1 U8373 ( .A(n4110), .B(\s13.dbus_out [53]), .C(n4109), .D(
        \s8.dbus_out [53]), .Z(n3907) );
  CND4X1 U8374 ( .A(n3910), .B(n3909), .C(n3908), .D(n3907), .Z(n1701) );
  CAOR2XL U8375 ( .A(\s1.addr [19]), .B(\s1.dbus_out [20]), .C(n4094), .D(
        \s7.dbus_out [20]), .Z(n3912) );
  CAOR2XL U8376 ( .A(\c1.Breset ), .B(data_stm_d[20]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [20]), .Z(n3911) );
  CANR3XL U8377 ( .A(\s6.addr [17]), .B(\s6.dbus_out [20]), .C(n3912), .D(
        n3911), .Z(n3921) );
  CND2X1 U8378 ( .A(n4098), .B(\s10.dbus_out [20]), .Z(n3916) );
  CANR2XL U8379 ( .A(n4078), .B(\s5.dbus_out [20]), .C(n4091), .D(
        \s4.dbus_out [20]), .Z(n3915) );
  CANR2XL U8380 ( .A(n4092), .B(\s14.dbus_out [20]), .C(\s12.dbus_out [20]), 
        .D(n4099), .Z(n3914) );
  CND2XL U8381 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [20]), .Z(n3913) );
  CAN4X1 U8382 ( .A(n3916), .B(n3915), .C(n3914), .D(n3913), .Z(n3920) );
  CAOR2XL U8383 ( .A(\s9.dbus_out [20]), .B(\s9.addr[16] ), .C(\s0.addr [14]), 
        .D(\s0.dbus_out [20]), .Z(n3917) );
  CANR1XL U8384 ( .A(n4108), .B(\s11.dbus_out [20]), .C(n3917), .Z(n3919) );
  CANR2X1 U8385 ( .A(n4110), .B(\s13.dbus_out [20]), .C(n4085), .D(
        \s8.dbus_out [20]), .Z(n3918) );
  CND4X1 U8386 ( .A(n3921), .B(n3920), .C(n3919), .D(n3918), .Z(n1734) );
  CAOR2XL U8387 ( .A(n4095), .B(\s1.dbus_out [21]), .C(n4094), .D(
        \s7.dbus_out [21]), .Z(n3923) );
  CAOR2XL U8388 ( .A(\c1.Breset ), .B(data_stm_d[21]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [21]), .Z(n3922) );
  CANR3X1 U8389 ( .A(\s6.addr [17]), .B(\s6.dbus_out [21]), .C(n3923), .D(
        n3922), .Z(n3933) );
  CNR2IX1 U8390 ( .B(\s10.dbus_out [21]), .A(n4076), .Z(n3924) );
  CIVX2 U8391 ( .A(n3924), .Z(n3928) );
  CANR2XL U8392 ( .A(n4078), .B(\s5.dbus_out [21]), .C(n4077), .D(
        \s4.dbus_out [21]), .Z(n3927) );
  CANR2XL U8393 ( .A(n4092), .B(\s14.dbus_out [21]), .C(\s12.dbus_out [21]), 
        .D(n4099), .Z(n3926) );
  CND2XL U8394 ( .A(n4101), .B(\s3.dbus_out [21]), .Z(n3925) );
  CAN4X1 U8395 ( .A(n3928), .B(n3927), .C(n3926), .D(n3925), .Z(n3932) );
  CAOR2XL U8396 ( .A(\s9.dbus_out [21]), .B(n5590), .C(n3940), .D(
        \s0.dbus_out [21]), .Z(n3929) );
  CANR1XL U8397 ( .A(n4093), .B(\s11.dbus_out [21]), .C(n3929), .Z(n3931) );
  CANR2XL U8398 ( .A(n4110), .B(\s13.dbus_out [21]), .C(\s8.en ), .D(
        \s8.dbus_out [21]), .Z(n3930) );
  CND4X1 U8399 ( .A(n3933), .B(n3932), .C(n3931), .D(n3930), .Z(n1733) );
  CAOR2XL U8400 ( .A(\s1.addr [19]), .B(\s1.dbus_out [22]), .C(n4094), .D(
        \s7.dbus_out [22]), .Z(n3935) );
  CAOR2XL U8401 ( .A(\c1.Breset ), .B(data_stm_d[22]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [22]), .Z(n3934) );
  CANR3X1 U8402 ( .A(n4075), .B(\s6.dbus_out [22]), .C(n3935), .D(n3934), .Z(
        n3945) );
  CANR2XL U8403 ( .A(n4078), .B(\s5.dbus_out [22]), .C(\s4.addr [19]), .D(
        \s4.dbus_out [22]), .Z(n3938) );
  CANR2XL U8404 ( .A(n4092), .B(\s14.dbus_out [22]), .C(\s12.dbus_out [22]), 
        .D(n4016), .Z(n3937) );
  CND2XL U8405 ( .A(n4101), .B(\s3.dbus_out [22]), .Z(n3936) );
  CAN4X1 U8406 ( .A(n3939), .B(n3938), .C(n3937), .D(n3936), .Z(n3944) );
  CAOR2XL U8407 ( .A(\s9.dbus_out [22]), .B(\s9.addr[8] ), .C(n3940), .D(
        \s0.dbus_out [22]), .Z(n3941) );
  CANR1XL U8408 ( .A(n4093), .B(\s11.dbus_out [22]), .C(n3941), .Z(n3943) );
  CANR2X1 U8409 ( .A(n4110), .B(\s13.dbus_out [22]), .C(n4109), .D(
        \s8.dbus_out [22]), .Z(n3942) );
  CND4X1 U8410 ( .A(n3945), .B(n3944), .C(n3943), .D(n3942), .Z(n1732) );
  CAOR2XL U8411 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [18]), .C(n4072), .D(
        \s7.dbus_out [18]), .Z(n3947) );
  CAOR2XL U8412 ( .A(\c1.Breset ), .B(data_stm_d[18]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [18]), .Z(n3946) );
  CANR3X1 U8413 ( .A(\s6.addr [17]), .B(\s6.dbus_out [18]), .C(n3947), .D(
        n3946), .Z(n3956) );
  CND2X1 U8414 ( .A(n4098), .B(\s10.dbus_out [18]), .Z(n3951) );
  CANR2XL U8415 ( .A(n4078), .B(\s5.dbus_out [18]), .C(n4077), .D(
        \s4.dbus_out [18]), .Z(n3950) );
  CANR2X1 U8416 ( .A(n4100), .B(\s14.dbus_out [18]), .C(\s12.dbus_out [18]), 
        .D(n4099), .Z(n3949) );
  CND2XL U8417 ( .A(n4101), .B(\s3.dbus_out [18]), .Z(n3948) );
  CAN4X1 U8418 ( .A(n3951), .B(n3950), .C(n3949), .D(n3948), .Z(n3955) );
  CAOR2XL U8419 ( .A(\s9.dbus_out [18]), .B(\s9.en ), .C(n3975), .D(
        \s0.dbus_out [18]), .Z(n3952) );
  CANR1XL U8420 ( .A(\s11.en ), .B(\s11.dbus_out [18]), .C(n3952), .Z(n3954)
         );
  CANR2X1 U8421 ( .A(n4110), .B(\s13.dbus_out [18]), .C(n4085), .D(
        \s8.dbus_out [18]), .Z(n3953) );
  CND4X1 U8422 ( .A(n3956), .B(n3955), .C(n3954), .D(n3953), .Z(n1736) );
  CAOR2X1 U8423 ( .A(n4090), .B(\s1.dbus_out [19]), .C(n4072), .D(
        \s7.dbus_out [19]), .Z(n3958) );
  CAOR2XL U8424 ( .A(\c1.Breset ), .B(data_stm_d[19]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [19]), .Z(n3957) );
  CANR3X1 U8425 ( .A(n1845), .B(\s6.dbus_out [19]), .C(n3958), .D(n3957), .Z(
        n3968) );
  CND2XL U8426 ( .A(\s10.en ), .B(\s10.dbus_out [19]), .Z(n3962) );
  CANR2XL U8427 ( .A(n4078), .B(\s5.dbus_out [19]), .C(n4077), .D(
        \s4.dbus_out [19]), .Z(n3961) );
  CANR2X1 U8428 ( .A(n4100), .B(\s14.dbus_out [19]), .C(\s12.dbus_out [19]), 
        .D(n4099), .Z(n3960) );
  CND2XL U8429 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [19]), .Z(n3959) );
  CAN4X1 U8430 ( .A(n3962), .B(n3961), .C(n3960), .D(n3959), .Z(n3967) );
  CAOR2XL U8431 ( .A(\s9.dbus_out [19]), .B(\s9.addr [15]), .C(n3963), .D(
        \s0.dbus_out [19]), .Z(n3964) );
  CANR1XL U8432 ( .A(n4093), .B(\s11.dbus_out [19]), .C(n3964), .Z(n3966) );
  CANR2X1 U8433 ( .A(n4110), .B(\s13.dbus_out [19]), .C(n4085), .D(
        \s8.dbus_out [19]), .Z(n3965) );
  CND4X1 U8434 ( .A(n3968), .B(n3967), .C(n3966), .D(n3965), .Z(n1735) );
  CAOR2XL U8435 ( .A(n4090), .B(\s1.dbus_out [24]), .C(\s7.en ), .D(
        \s7.dbus_out [24]), .Z(n3970) );
  CAOR2XL U8436 ( .A(\c1.Breset ), .B(data_stm_d[24]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [24]), .Z(n3969) );
  CANR3X1 U8437 ( .A(n1845), .B(\s6.dbus_out [24]), .C(n3970), .D(n3969), .Z(
        n3980) );
  CND2X1 U8438 ( .A(n4098), .B(\s10.dbus_out [24]), .Z(n3974) );
  CANR2XL U8439 ( .A(n4078), .B(\s5.dbus_out [24]), .C(n4091), .D(
        \s4.dbus_out [24]), .Z(n3973) );
  CANR2XL U8440 ( .A(n4100), .B(\s14.dbus_out [24]), .C(\s12.dbus_out [24]), 
        .D(n4099), .Z(n3972) );
  CND2XL U8441 ( .A(\s3.addr [18]), .B(\s3.dbus_out [24]), .Z(n3971) );
  CAN4X1 U8442 ( .A(n3974), .B(n3973), .C(n3972), .D(n3971), .Z(n3979) );
  CAOR2XL U8443 ( .A(\s9.dbus_out [24]), .B(\s9.addr[7] ), .C(n3975), .D(
        \s0.dbus_out [24]), .Z(n3976) );
  CANR1XL U8444 ( .A(n4093), .B(\s11.dbus_out [24]), .C(n3976), .Z(n3978) );
  CANR2X1 U8445 ( .A(n4110), .B(\s13.dbus_out [24]), .C(n4085), .D(
        \s8.dbus_out [24]), .Z(n3977) );
  CND4X1 U8446 ( .A(n3980), .B(n3979), .C(n3978), .D(n3977), .Z(n1730) );
  CAOR2XL U8447 ( .A(n4090), .B(\s1.dbus_out [25]), .C(n4072), .D(
        \s7.dbus_out [25]), .Z(n3982) );
  CAOR2XL U8448 ( .A(\c1.Breset ), .B(data_stm_d[25]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [25]), .Z(n3981) );
  CANR3X1 U8449 ( .A(n1845), .B(\s6.dbus_out [25]), .C(n3982), .D(n3981), .Z(
        n3991) );
  CND2XL U8450 ( .A(\s10.en ), .B(\s10.dbus_out [25]), .Z(n3986) );
  CANR2XL U8451 ( .A(n4078), .B(\s5.dbus_out [25]), .C(n4077), .D(
        \s4.dbus_out [25]), .Z(n3985) );
  CANR2X1 U8452 ( .A(n4092), .B(\s14.dbus_out [25]), .C(\s12.dbus_out [25]), 
        .D(n4099), .Z(n3984) );
  CND2XL U8453 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [25]), .Z(n3983) );
  CAN4X1 U8454 ( .A(n3986), .B(n3985), .C(n3984), .D(n3983), .Z(n3990) );
  CAOR2XL U8455 ( .A(\s9.dbus_out [25]), .B(\s9.addr[16] ), .C(\s0.addr [13]), 
        .D(\s0.dbus_out [25]), .Z(n3987) );
  CANR1XL U8456 ( .A(n4093), .B(\s11.dbus_out [25]), .C(n3987), .Z(n3989) );
  CANR2X1 U8457 ( .A(n4110), .B(\s13.dbus_out [25]), .C(n4109), .D(
        \s8.dbus_out [25]), .Z(n3988) );
  CND4X1 U8458 ( .A(n3991), .B(n3990), .C(n3989), .D(n3988), .Z(n1729) );
  CAOR2XL U8459 ( .A(n4090), .B(\s1.dbus_out [32]), .C(n4094), .D(
        \s7.dbus_out [32]), .Z(n3993) );
  CAOR2XL U8460 ( .A(\c1.Breset ), .B(data_stm_d[32]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [32]), .Z(n3992) );
  CANR3X1 U8461 ( .A(n4075), .B(\s6.dbus_out [32]), .C(n3993), .D(n3992), .Z(
        n4002) );
  CND2X1 U8462 ( .A(n4098), .B(\s10.dbus_out [32]), .Z(n3997) );
  CANR2X1 U8463 ( .A(n4078), .B(\s5.dbus_out [32]), .C(n4091), .D(
        \s4.dbus_out [32]), .Z(n3996) );
  CANR2X1 U8464 ( .A(n4092), .B(\s14.dbus_out [32]), .C(\s12.dbus_out [32]), 
        .D(n4099), .Z(n3995) );
  CND2XL U8465 ( .A(\s3.addr[14] ), .B(\s3.dbus_out [32]), .Z(n3994) );
  CAN4X1 U8466 ( .A(n3997), .B(n3996), .C(n3995), .D(n3994), .Z(n4001) );
  CAOR2XL U8467 ( .A(\s9.dbus_out [32]), .B(\s9.addr[8] ), .C(\s0.en ), .D(
        \s0.dbus_out [32]), .Z(n3998) );
  CANR1XL U8468 ( .A(n4093), .B(\s11.dbus_out [32]), .C(n3998), .Z(n4000) );
  CANR2XL U8469 ( .A(n4110), .B(\s13.dbus_out [32]), .C(n4109), .D(
        \s8.dbus_out [32]), .Z(n3999) );
  CND4X1 U8470 ( .A(n4002), .B(n4001), .C(n4000), .D(n3999), .Z(n1722) );
  CAOR2XL U8471 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [27]), .C(n4094), .D(
        \s7.dbus_out [27]), .Z(n4004) );
  CAOR2XL U8472 ( .A(\c1.Breset ), .B(data_stm_d[27]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [27]), .Z(n4003) );
  CANR3X1 U8473 ( .A(n1845), .B(\s6.dbus_out [27]), .C(n4004), .D(n4003), .Z(
        n4013) );
  CND2XL U8474 ( .A(n4098), .B(\s10.dbus_out [27]), .Z(n4008) );
  CANR2X1 U8475 ( .A(n4078), .B(\s5.dbus_out [27]), .C(n4077), .D(
        \s4.dbus_out [27]), .Z(n4007) );
  CANR2XL U8476 ( .A(n4092), .B(\s14.dbus_out [27]), .C(\s12.dbus_out [27]), 
        .D(n1843), .Z(n4006) );
  CND2XL U8477 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [27]), .Z(n4005) );
  CAN4X1 U8478 ( .A(n4008), .B(n4007), .C(n4006), .D(n4005), .Z(n4012) );
  CAOR2XL U8479 ( .A(\s9.dbus_out [27]), .B(\s9.addr[7] ), .C(\s0.addr [14]), 
        .D(\s0.dbus_out [27]), .Z(n4009) );
  CANR1XL U8480 ( .A(n4093), .B(\s11.dbus_out [27]), .C(n4009), .Z(n4011) );
  CANR2X1 U8481 ( .A(n4110), .B(\s13.dbus_out [27]), .C(n4109), .D(
        \s8.dbus_out [27]), .Z(n4010) );
  CND4X1 U8482 ( .A(n4013), .B(n4012), .C(n4011), .D(n4010), .Z(n1727) );
  CAOR2X1 U8483 ( .A(n4095), .B(\s1.dbus_out [41]), .C(n4072), .D(
        \s7.dbus_out [41]), .Z(n4015) );
  CAOR2XL U8484 ( .A(\c1.Breset ), .B(data_stm_d[41]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [41]), .Z(n4014) );
  CANR3X1 U8485 ( .A(n1845), .B(\s6.dbus_out [41]), .C(n4015), .D(n4014), .Z(
        n4025) );
  CANR2XL U8486 ( .A(n4078), .B(\s5.dbus_out [41]), .C(n4077), .D(
        \s4.dbus_out [41]), .Z(n4019) );
  CANR2XL U8487 ( .A(n4100), .B(\s14.dbus_out [41]), .C(\s12.dbus_out [41]), 
        .D(n4016), .Z(n4018) );
  CND2X1 U8488 ( .A(n4101), .B(\s3.dbus_out [41]), .Z(n4017) );
  CAN4X1 U8489 ( .A(n4020), .B(n4019), .C(n4018), .D(n4017), .Z(n4024) );
  CAOR2XL U8490 ( .A(\s9.dbus_out [41]), .B(\s9.addr[8] ), .C(\s0.addr [14]), 
        .D(\s0.dbus_out [41]), .Z(n4021) );
  CANR1XL U8491 ( .A(n4108), .B(\s11.dbus_out [41]), .C(n4021), .Z(n4023) );
  CANR2X1 U8492 ( .A(n4110), .B(\s13.dbus_out [41]), .C(n4109), .D(
        \s8.dbus_out [41]), .Z(n4022) );
  CND4X1 U8493 ( .A(n4025), .B(n4024), .C(n4023), .D(n4022), .Z(n1713) );
  CAOR2X1 U8494 ( .A(n4090), .B(\s1.dbus_out [34]), .C(n4094), .D(
        \s7.dbus_out [34]), .Z(n4027) );
  CAOR2XL U8495 ( .A(\c1.Breset ), .B(data_stm_d[34]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [34]), .Z(n4026) );
  CANR3XL U8496 ( .A(n4062), .B(\s6.dbus_out [34]), .C(n4027), .D(n4026), .Z(
        n4036) );
  CND2XL U8497 ( .A(\s10.en ), .B(\s10.dbus_out [34]), .Z(n4031) );
  CANR2XL U8498 ( .A(n4078), .B(\s5.dbus_out [34]), .C(n4077), .D(
        \s4.dbus_out [34]), .Z(n4030) );
  CANR2X1 U8499 ( .A(n4092), .B(\s14.dbus_out [34]), .C(\s12.dbus_out [34]), 
        .D(n4099), .Z(n4029) );
  CND2XL U8500 ( .A(\s3.addr [18]), .B(\s3.dbus_out [34]), .Z(n4028) );
  CAN4X1 U8501 ( .A(n4031), .B(n4030), .C(n4029), .D(n4028), .Z(n4035) );
  CAOR2XL U8502 ( .A(\s9.dbus_out [34]), .B(\s9.addr [15]), .C(\s0.addr [12]), 
        .D(\s0.dbus_out [34]), .Z(n4032) );
  CANR1XL U8503 ( .A(\s11.dbus_out [34]), .B(\s11.addr[17] ), .C(n4032), .Z(
        n4034) );
  CANR2XL U8504 ( .A(n4110), .B(\s13.dbus_out [34]), .C(\s8.en ), .D(
        \s8.dbus_out [34]), .Z(n4033) );
  CND4X1 U8505 ( .A(n4036), .B(n4035), .C(n4034), .D(n4033), .Z(n1720) );
  CAOR2XL U8506 ( .A(n4090), .B(\s1.dbus_out [42]), .C(n4094), .D(
        \s7.dbus_out [42]), .Z(n4038) );
  CAOR2XL U8507 ( .A(\c1.Breset ), .B(data_stm_d[42]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [42]), .Z(n4037) );
  CANR3X1 U8508 ( .A(n1845), .B(\s6.dbus_out [42]), .C(n4038), .D(n4037), .Z(
        n4047) );
  CND2XL U8509 ( .A(\s10.en ), .B(\s10.dbus_out [42]), .Z(n4042) );
  CANR2X1 U8510 ( .A(n4078), .B(\s5.dbus_out [42]), .C(n4077), .D(
        \s4.dbus_out [42]), .Z(n4041) );
  CANR2XL U8511 ( .A(n4100), .B(\s14.dbus_out [42]), .C(\s12.dbus_out [42]), 
        .D(n1843), .Z(n4040) );
  CND2XL U8512 ( .A(\s3.addr [18]), .B(\s3.dbus_out [42]), .Z(n4039) );
  CAN4X1 U8513 ( .A(n4042), .B(n4041), .C(n4040), .D(n4039), .Z(n4046) );
  CAOR2XL U8514 ( .A(\s9.dbus_out [42]), .B(\s9.addr[8] ), .C(\s0.addr [12]), 
        .D(\s0.dbus_out [42]), .Z(n4043) );
  CANR1XL U8515 ( .A(n4093), .B(\s11.dbus_out [42]), .C(n4043), .Z(n4045) );
  CANR2XL U8516 ( .A(n4110), .B(\s13.dbus_out [42]), .C(\s8.dbus_out [42]), 
        .D(n4085), .Z(n4044) );
  CND4X1 U8517 ( .A(n4047), .B(n4046), .C(n4045), .D(n4044), .Z(n1712) );
  CAOR2XL U8518 ( .A(\s1.addr [19]), .B(\s1.dbus_out [28]), .C(n4072), .D(
        \s7.dbus_out [28]), .Z(n4049) );
  CAOR2XL U8519 ( .A(\c1.Breset ), .B(data_stm_d[28]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [28]), .Z(n4048) );
  CANR3X1 U8520 ( .A(n4075), .B(\s6.dbus_out [28]), .C(n4049), .D(n4048), .Z(
        n4059) );
  CND2XL U8521 ( .A(n4098), .B(\s10.dbus_out [28]), .Z(n4054) );
  CANR2XL U8522 ( .A(n4078), .B(\s5.dbus_out [28]), .C(n4077), .D(
        \s4.dbus_out [28]), .Z(n4053) );
  CANR2XL U8523 ( .A(\s14.addr[16] ), .B(\s14.dbus_out [28]), .C(
        \s12.dbus_out [28]), .D(n4099), .Z(n4052) );
  CND2XL U8524 ( .A(\s3.addr[9] ), .B(\s3.dbus_out [28]), .Z(n4051) );
  CAN4X1 U8525 ( .A(n4054), .B(n4053), .C(n4052), .D(n4051), .Z(n4058) );
  CAOR2XL U8526 ( .A(\s9.dbus_out [28]), .B(\s9.en ), .C(\s0.addr [13]), .D(
        \s0.dbus_out [28]), .Z(n4055) );
  CANR1XL U8527 ( .A(n4108), .B(\s11.dbus_out [28]), .C(n4055), .Z(n4057) );
  CANR2X1 U8528 ( .A(n4110), .B(\s13.dbus_out [28]), .C(n4085), .D(
        \s8.dbus_out [28]), .Z(n4056) );
  CND4X1 U8529 ( .A(n4059), .B(n4058), .C(n4057), .D(n4056), .Z(n1726) );
  CAOR2XL U8530 ( .A(\s1.addr[17] ), .B(\s1.dbus_out [43]), .C(n4094), .D(
        \s7.dbus_out [43]), .Z(n4061) );
  CAOR2XL U8531 ( .A(\c1.Breset ), .B(data_stm_d[43]), .C(\s2.addr[16] ), .D(
        \s2.dbus_out [43]), .Z(n4060) );
  CANR3XL U8532 ( .A(n4062), .B(\s6.dbus_out [43]), .C(n4061), .D(n4060), .Z(
        n4071) );
  CND2X1 U8533 ( .A(n4098), .B(\s10.dbus_out [43]), .Z(n4066) );
  CANR2XL U8534 ( .A(n4078), .B(\s5.dbus_out [43]), .C(n4091), .D(
        \s4.dbus_out [43]), .Z(n4065) );
  CANR2XL U8535 ( .A(n4100), .B(\s14.dbus_out [43]), .C(\s12.dbus_out [43]), 
        .D(n4099), .Z(n4064) );
  CND2XL U8536 ( .A(n4101), .B(\s3.dbus_out [43]), .Z(n4063) );
  CAN4X1 U8537 ( .A(n4066), .B(n4065), .C(n4064), .D(n4063), .Z(n4070) );
  CAOR2XL U8538 ( .A(\s9.dbus_out [43]), .B(\s9.addr[7] ), .C(n4083), .D(
        \s0.dbus_out [43]), .Z(n4067) );
  CANR1XL U8539 ( .A(n4093), .B(\s11.dbus_out [43]), .C(n4067), .Z(n4069) );
  CANR2XL U8540 ( .A(n4110), .B(\s13.dbus_out [43]), .C(\s8.en ), .D(
        \s8.dbus_out [43]), .Z(n4068) );
  CND4X1 U8541 ( .A(n4071), .B(n4070), .C(n4069), .D(n4068), .Z(n1711) );
  CAOR2XL U8542 ( .A(\s1.addr [19]), .B(\s1.dbus_out [29]), .C(n4072), .D(
        \s7.dbus_out [29]), .Z(n4074) );
  CAOR2XL U8543 ( .A(\c1.Breset ), .B(data_stm_d[29]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [29]), .Z(n4073) );
  CANR3X1 U8544 ( .A(n4075), .B(\s6.dbus_out [29]), .C(n4074), .D(n4073), .Z(
        n4089) );
  CANR2XL U8545 ( .A(n4078), .B(\s5.dbus_out [29]), .C(n4077), .D(
        \s4.dbus_out [29]), .Z(n4081) );
  CANR2X1 U8546 ( .A(n4100), .B(\s14.dbus_out [29]), .C(\s12.dbus_out [29]), 
        .D(n4099), .Z(n4080) );
  CND2XL U8547 ( .A(n4101), .B(\s3.dbus_out [29]), .Z(n4079) );
  CAN4X1 U8548 ( .A(n4082), .B(n4081), .C(n4080), .D(n4079), .Z(n4088) );
  CAOR2XL U8549 ( .A(\s9.dbus_out [29]), .B(\s9.addr[7] ), .C(n4083), .D(
        \s0.dbus_out [29]), .Z(n4084) );
  CANR1XL U8550 ( .A(n4093), .B(\s11.dbus_out [29]), .C(n4084), .Z(n4087) );
  CANR2XL U8551 ( .A(n4110), .B(\s13.dbus_out [29]), .C(n4085), .D(
        \s8.dbus_out [29]), .Z(n4086) );
  CND4X1 U8552 ( .A(n4089), .B(n4088), .C(n4087), .D(n4086), .Z(n1725) );
  CAOR2XL U8553 ( .A(n4095), .B(\s1.dbus_out [23]), .C(n4094), .D(
        \s7.dbus_out [23]), .Z(n4097) );
  CAOR2XL U8554 ( .A(\c1.Breset ), .B(data_stm_d[23]), .C(\s2.addr[19] ), .D(
        \s2.dbus_out [23]), .Z(n4096) );
  CANR3X1 U8555 ( .A(n1845), .B(\s6.dbus_out [23]), .C(n4097), .D(n4096), .Z(
        n4114) );
  CND2X1 U8556 ( .A(n4098), .B(\s10.dbus_out [23]), .Z(n4105) );
  CANR2XL U8557 ( .A(n4078), .B(\s5.dbus_out [23]), .C(\s4.addr [19]), .D(
        \s4.dbus_out [23]), .Z(n4104) );
  CANR2XL U8558 ( .A(n4100), .B(\s14.dbus_out [23]), .C(\s12.dbus_out [23]), 
        .D(n4099), .Z(n4103) );
  CND2XL U8559 ( .A(n4101), .B(\s3.dbus_out [23]), .Z(n4102) );
  CAN4X1 U8560 ( .A(n4105), .B(n4104), .C(n4103), .D(n4102), .Z(n4113) );
  CAOR2XL U8561 ( .A(\s9.dbus_out [23]), .B(\s9.addr[7] ), .C(n4106), .D(
        \s0.dbus_out [23]), .Z(n4107) );
  CANR1XL U8562 ( .A(n4108), .B(\s11.dbus_out [23]), .C(n4107), .Z(n4112) );
  CANR2X1 U8563 ( .A(n4110), .B(\s13.dbus_out [23]), .C(n4109), .D(
        \s8.dbus_out [23]), .Z(n4111) );
  CND4X1 U8564 ( .A(n4114), .B(n4113), .C(n4112), .D(n4111), .Z(n1731) );
  CIVX2 U8565 ( .A(n4115), .Z(n4183) );
  CNR2X1 U8566 ( .A(n4255), .B(n4183), .Z(\s2.SbusIn [10]) );
  CIVX2 U8567 ( .A(n4116), .Z(n4316) );
  CNR2X1 U8568 ( .A(n4255), .B(n4316), .Z(\s2.SbusIn [8]) );
  CIVX2 U8569 ( .A(n4117), .Z(n4273) );
  CNR2X1 U8570 ( .A(n4255), .B(n4273), .Z(\s2.SbusIn [28]) );
  CIVX2 U8571 ( .A(n4118), .Z(n4206) );
  CNR2X1 U8572 ( .A(n4255), .B(n4206), .Z(\s2.addr [23]) );
  CIVX2 U8573 ( .A(n4119), .Z(n4292) );
  CNR2X1 U8574 ( .A(n4255), .B(n4292), .Z(\s2.SbusIn [31]) );
  CIVX2 U8575 ( .A(n4120), .Z(n4261) );
  CNR2X1 U8576 ( .A(n4256), .B(n4261), .Z(\s2.SbusIn [63]) );
  CIVX2 U8577 ( .A(n4121), .Z(n4226) );
  CNR2X1 U8578 ( .A(n4256), .B(n4226), .Z(\s2.SbusIn [48]) );
  CIVX2 U8579 ( .A(n4122), .Z(n4284) );
  CNR2X1 U8580 ( .A(n4256), .B(n4284), .Z(\s2.addr [43]) );
  CIVX2 U8581 ( .A(n4123), .Z(n4247) );
  CNR2X1 U8582 ( .A(n4256), .B(n4247), .Z(\s2.SbusIn [13]) );
  CIVX2 U8583 ( .A(n4124), .Z(n4322) );
  CNR2X1 U8584 ( .A(n4256), .B(n4322), .Z(\s2.addr [36]) );
  CIVX2 U8585 ( .A(n4125), .Z(n4191) );
  CNR2X1 U8586 ( .A(n4255), .B(n4191), .Z(\s2.SbusIn [61]) );
  CNR2X1 U8587 ( .A(n4255), .B(n4289), .Z(\s2.SbusIn [46]) );
  CIVX2 U8588 ( .A(n4126), .Z(n4211) );
  CNR2X1 U8589 ( .A(n4255), .B(n4211), .Z(\s2.SbusIn [62]) );
  CIVX2 U8590 ( .A(n4127), .Z(n4249) );
  CNR2X1 U8591 ( .A(n4255), .B(n4249), .Z(\s2.SbusIn [50]) );
  CIVX2 U8592 ( .A(n4128), .Z(n4184) );
  CNR2X1 U8593 ( .A(n4256), .B(n4184), .Z(\s2.addr [21]) );
  CIVX2 U8594 ( .A(n4129), .Z(n4303) );
  CNR2X1 U8595 ( .A(n4255), .B(n4303), .Z(\s2.SbusIn [45]) );
  CIVX2 U8596 ( .A(n4130), .Z(n4219) );
  CNR2X1 U8597 ( .A(n4256), .B(n4219), .Z(\s2.SbusIn [59]) );
  CIVX2 U8598 ( .A(n4131), .Z(n4221) );
  CNR2X1 U8599 ( .A(n4256), .B(n4221), .Z(\s2.addr [34]) );
  CIVX2 U8600 ( .A(n4132), .Z(n4286) );
  CNR2X1 U8601 ( .A(n4255), .B(n4286), .Z(\s2.SbusIn [43]) );
  CNR2X1 U8602 ( .A(n4256), .B(n4312), .Z(\s2.addr [40]) );
  CIVX2 U8603 ( .A(n4133), .Z(n4217) );
  CNR2X1 U8604 ( .A(n4255), .B(n4217), .Z(\s2.addr [28]) );
  CIVX2 U8605 ( .A(n4134), .Z(n4182) );
  CNR2X1 U8606 ( .A(n4255), .B(n4182), .Z(\s2.addr [29]) );
  CIVX2 U8607 ( .A(n4135), .Z(n4293) );
  CNR2X1 U8608 ( .A(n4256), .B(n4293), .Z(\s2.SbusIn [39]) );
  CIVX2 U8609 ( .A(n4136), .Z(n4189) );
  CNR2X1 U8610 ( .A(n4256), .B(n4189), .Z(\s2.addr [46]) );
  CIVX2 U8611 ( .A(n4331), .Z(n4205) );
  CNR2X1 U8612 ( .A(n4255), .B(n4205), .Z(\s2.addr [20]) );
  CIVX2 U8613 ( .A(n4137), .Z(n4203) );
  CNR2X1 U8614 ( .A(n4256), .B(n4203), .Z(\s2.addr [48]) );
  CNR2X1 U8615 ( .A(n4256), .B(n4230), .Z(\s2.addr [22]) );
  CIVX2 U8616 ( .A(n4138), .Z(n4320) );
  CNR2X1 U8617 ( .A(n4256), .B(n4320), .Z(\s2.SbusIn [44]) );
  CIVX2 U8618 ( .A(n4139), .Z(n4218) );
  CNR2X1 U8619 ( .A(n4255), .B(n4218), .Z(\s2.SbusIn [47]) );
  CNR2X1 U8620 ( .A(n4255), .B(n4250), .Z(\s2.addr [62]) );
  CIVX2 U8621 ( .A(n4140), .Z(n4229) );
  CNR2X1 U8622 ( .A(n4256), .B(n4229), .Z(\s2.addr [63]) );
  CIVX2 U8623 ( .A(n4141), .Z(n4181) );
  CNR2X1 U8624 ( .A(n4255), .B(n4181), .Z(\s2.SbusIn [25]) );
  CNR2X1 U8625 ( .A(n4255), .B(n4302), .Z(\s2.SbusIn [12]) );
  CNR2X1 U8626 ( .A(n4255), .B(n4210), .Z(\s2.SbusIn [23]) );
  CNR2X1 U8627 ( .A(n4256), .B(n4209), .Z(\s2.SbusIn [11]) );
  CNR2X1 U8628 ( .A(n4256), .B(n4257), .Z(\s2.addr [7]) );
  CIVX2 U8629 ( .A(n4142), .Z(n4269) );
  CNR2X1 U8630 ( .A(n4256), .B(n4269), .Z(\s2.SbusIn [41]) );
  CNR2X1 U8631 ( .A(n4255), .B(n4300), .Z(\s2.addr [41]) );
  CIVX2 U8632 ( .A(n4143), .Z(n4265) );
  CNR2X1 U8633 ( .A(n4255), .B(n4265), .Z(\s2.SbusIn [40]) );
  CIVX2 U8634 ( .A(n4144), .Z(n4299) );
  CNR2X1 U8635 ( .A(n4255), .B(n4299), .Z(\s2.SbusIn [42]) );
  CIVX2 U8636 ( .A(n4145), .Z(n4304) );
  CNR2X1 U8637 ( .A(n4256), .B(n4304), .Z(\s2.SbusIn [30]) );
  CIVX2 U8638 ( .A(n4146), .Z(n4186) );
  CNR2X1 U8639 ( .A(n4256), .B(n4186), .Z(\s2.addr [47]) );
  CNR2X1 U8640 ( .A(n4256), .B(n4212), .Z(\s2.SbusIn [27]) );
  CIVX2 U8641 ( .A(n4147), .Z(n4248) );
  CNR2X1 U8642 ( .A(n4256), .B(n4248), .Z(\s2.SbusIn [26]) );
  CIVX2 U8643 ( .A(n4148), .Z(n4252) );
  CNR2X1 U8644 ( .A(n4255), .B(n4252), .Z(\s2.addr [54]) );
  CIVX2 U8645 ( .A(n4149), .Z(n4280) );
  CNR2X1 U8646 ( .A(n4256), .B(n4280), .Z(\s2.SbusIn [24]) );
  CNR2X1 U8647 ( .A(n4256), .B(n4228), .Z(\s2.SbusIn [5]) );
  CIVX2 U8648 ( .A(n4150), .Z(n4295) );
  CNR2X1 U8649 ( .A(n4255), .B(n4295), .Z(\s2.SbusIn [20]) );
  CIVX2 U8650 ( .A(n4151), .Z(n4296) );
  CNR2X1 U8651 ( .A(n4255), .B(n4296), .Z(\s2.addr [61]) );
  CIVX2 U8652 ( .A(n4152), .Z(n4222) );
  CNR2X1 U8653 ( .A(n4255), .B(n4222), .Z(\s2.SbusIn [19]) );
  CIVX2 U8654 ( .A(n4329), .Z(n4187) );
  CNR2X1 U8655 ( .A(n4255), .B(n4187), .Z(\s2.SbusIn [6]) );
  CIVX2 U8656 ( .A(n4153), .Z(n4223) );
  CNR2X1 U8657 ( .A(n4255), .B(n4223), .Z(\s2.addr [42]) );
  CIVX2 U8658 ( .A(n4154), .Z(n4268) );
  CNR2X1 U8659 ( .A(n4256), .B(n4268), .Z(\s2.SbusIn [7]) );
  CIVX2 U8660 ( .A(n4155), .Z(n4275) );
  CNR2X1 U8661 ( .A(n4256), .B(n4275), .Z(\s2.addr [49]) );
  CIVX2 U8662 ( .A(n4156), .Z(n4240) );
  CNR2X1 U8663 ( .A(n4258), .B(n4240), .Z(\s13.SbusIn [33]) );
  CNR2X1 U8664 ( .A(n4258), .B(n4187), .Z(\s13.SbusIn [6]) );
  CNR2X1 U8665 ( .A(n4259), .B(n4322), .Z(\s13.addr [36]) );
  CNR2X1 U8666 ( .A(n4259), .B(n4318), .Z(\s13.addr [2]) );
  CIVX2 U8667 ( .A(n4157), .Z(n4287) );
  CNR2X1 U8668 ( .A(n4258), .B(n4287), .Z(\s13.addr [32]) );
  CNR2X1 U8669 ( .A(n4258), .B(n4303), .Z(\s13.SbusIn [45]) );
  CIVX2 U8670 ( .A(n4158), .Z(n4227) );
  CNR2X1 U8671 ( .A(n4259), .B(n4227), .Z(\s13.SbusIn [21]) );
  CNR2X1 U8672 ( .A(n4259), .B(n4226), .Z(\s13.SbusIn [48]) );
  CIVX2 U8673 ( .A(n4159), .Z(n4283) );
  CNR2X1 U8674 ( .A(n4258), .B(n4283), .Z(\s13.SbusIn [56]) );
  CIVX2 U8675 ( .A(n4160), .Z(n4305) );
  CNR2X1 U8676 ( .A(n4258), .B(n4305), .Z(\s13.addr [31]) );
  CNR2X1 U8677 ( .A(n4259), .B(n4261), .Z(\s13.SbusIn [63]) );
  CNR2X1 U8678 ( .A(n4258), .B(n4221), .Z(\s13.addr [34]) );
  CNR2X1 U8679 ( .A(n4259), .B(n4191), .Z(\s13.SbusIn [61]) );
  CNR2X1 U8680 ( .A(n4259), .B(n4182), .Z(\s13.addr [29]) );
  CNR2X1 U8681 ( .A(n4258), .B(n4223), .Z(\s13.addr [42]) );
  CIVX2 U8682 ( .A(n4161), .Z(n4294) );
  CNR2X1 U8683 ( .A(n4259), .B(n4294), .Z(\s13.SbusIn [57]) );
  CNR2X1 U8684 ( .A(n4259), .B(n4284), .Z(\s13.addr [43]) );
  CNR2X1 U8685 ( .A(n4258), .B(n4324), .Z(\s13.addr [44]) );
  CIVX2 U8686 ( .A(n4162), .Z(n4238) );
  CNR2X1 U8687 ( .A(n4258), .B(n4238), .Z(\s13.addr [45]) );
  CNR2X1 U8688 ( .A(n4258), .B(n4189), .Z(\s13.addr [46]) );
  CIVX2 U8689 ( .A(n4163), .Z(n4233) );
  CNR2X1 U8690 ( .A(n4259), .B(n4233), .Z(\s13.SbusIn [51]) );
  CNR2X1 U8691 ( .A(n4258), .B(n4186), .Z(\s13.addr [47]) );
  CNR2X1 U8692 ( .A(n4259), .B(n4203), .Z(\s13.addr [48]) );
  CNR2X1 U8693 ( .A(n4259), .B(n4217), .Z(\s13.addr [28]) );
  CIVX2 U8694 ( .A(n4164), .Z(n4260) );
  CNR2X1 U8695 ( .A(n4258), .B(n4260), .Z(\s13.addr [50]) );
  CIVX2 U8696 ( .A(n4165), .Z(n4264) );
  CNR2X1 U8697 ( .A(n4259), .B(n4264), .Z(\s13.addr [51]) );
  CIVX2 U8698 ( .A(n4166), .Z(n4276) );
  CNR2X1 U8699 ( .A(n4258), .B(n4276), .Z(\s13.addr [52]) );
  CNR2X1 U8700 ( .A(n4259), .B(n4269), .Z(\s13.SbusIn [41]) );
  CNR2X1 U8701 ( .A(n4258), .B(n4299), .Z(\s13.SbusIn [42]) );
  CNR2X1 U8702 ( .A(n4259), .B(n4209), .Z(\s13.SbusIn [11]) );
  CNR2X1 U8703 ( .A(n4258), .B(n4272), .Z(\s13.addr [0]) );
  CNR2X1 U8704 ( .A(n4259), .B(n4212), .Z(\s13.SbusIn [27]) );
  CNR2X1 U8705 ( .A(n4259), .B(n4181), .Z(\s13.SbusIn [25]) );
  CNR2X1 U8706 ( .A(n4258), .B(n4273), .Z(\s13.SbusIn [28]) );
  CNR2X1 U8707 ( .A(n4259), .B(n4288), .Z(\s13.SbusIn [16]) );
  CNR2X1 U8708 ( .A(n4258), .B(n4211), .Z(\s13.SbusIn [62]) );
  CNR2X1 U8709 ( .A(n4259), .B(n4225), .Z(\s13.SbusIn [14]) );
  CIVX2 U8710 ( .A(n4167), .Z(n4235) );
  CNR2X1 U8711 ( .A(n4259), .B(n4235), .Z(\s13.SbusIn [60]) );
  CIVX2 U8712 ( .A(n4168), .Z(n4234) );
  CNR2X1 U8713 ( .A(n4258), .B(n4234), .Z(\s13.SbusIn [58]) );
  CNR2X1 U8714 ( .A(n4258), .B(n4286), .Z(\s13.SbusIn [43]) );
  CIVX2 U8715 ( .A(n4169), .Z(n4297) );
  CNR2X1 U8716 ( .A(n4259), .B(n4297), .Z(\s13.SbusIn [15]) );
  CNR2X1 U8717 ( .A(n4258), .B(n4265), .Z(\s13.SbusIn [40]) );
  CIVX2 U8718 ( .A(n4170), .Z(n4271) );
  CNR2X1 U8719 ( .A(n4258), .B(n4271), .Z(\s13.SbusIn [53]) );
  CNR2X1 U8720 ( .A(n4259), .B(n4213), .Z(\s13.SbusIn [52]) );
  CNR2X1 U8721 ( .A(n4258), .B(n4183), .Z(\s13.SbusIn [10]) );
  CIVX2 U8722 ( .A(n4171), .Z(n4298) );
  CNR2X1 U8723 ( .A(n4258), .B(n4298), .Z(\s13.SbusIn [32]) );
  CNR2X1 U8724 ( .A(n4258), .B(n4218), .Z(\s13.SbusIn [47]) );
  CNR2X1 U8725 ( .A(n4259), .B(n4320), .Z(\s13.SbusIn [44]) );
  CIVX2 U8726 ( .A(n4172), .Z(n4310) );
  CNR2X1 U8727 ( .A(n4259), .B(n4310), .Z(\s13.SbusIn [17]) );
  CIVX2 U8728 ( .A(n4173), .Z(n4216) );
  CNR2X1 U8729 ( .A(n4258), .B(n4216), .Z(\s13.addr [35]) );
  CIVX2 U8730 ( .A(n4174), .Z(n4239) );
  CNR2X1 U8731 ( .A(n4258), .B(n4239), .Z(\s13.addr [53]) );
  CIVX2 U8732 ( .A(n4175), .Z(n4263) );
  CNR2X1 U8733 ( .A(n4259), .B(n4263), .Z(\s13.SbusIn [54]) );
  CNR2X1 U8734 ( .A(n4259), .B(n4228), .Z(\s13.SbusIn [5]) );
  CNR2X1 U8735 ( .A(n4258), .B(n4308), .Z(\s13.SbusIn [55]) );
  CIVX2 U8736 ( .A(n4176), .Z(n4236) );
  CNR2X1 U8737 ( .A(n4258), .B(n4236), .Z(\s13.addr [30]) );
  CNR2X1 U8738 ( .A(n4259), .B(n4184), .Z(\s13.addr [21]) );
  CNR2X1 U8739 ( .A(n4259), .B(n4205), .Z(\s13.addr [20]) );
  CNR2X1 U8740 ( .A(n4258), .B(n4312), .Z(\s13.addr [40]) );
  CNR2X1 U8741 ( .A(n4259), .B(n4289), .Z(\s13.SbusIn [46]) );
  CIVX2 U8742 ( .A(n4177), .Z(n4267) );
  CNR2X1 U8743 ( .A(n4259), .B(n4267), .Z(\s13.addr [39]) );
  CNR2X1 U8744 ( .A(n4258), .B(n4285), .Z(\s13.addr [37]) );
  CIVX2 U8745 ( .A(n4178), .Z(n4220) );
  CNR2X1 U8746 ( .A(n4258), .B(n4220), .Z(\s13.SbusIn [34]) );
  CNR2X1 U8747 ( .A(n4259), .B(n4304), .Z(\s13.SbusIn [30]) );
  CIVX2 U8748 ( .A(n4179), .Z(n4306) );
  CNR2X1 U8749 ( .A(n4259), .B(n4306), .Z(\s13.addr [33]) );
  CNR2X1 U8750 ( .A(n4258), .B(n4231), .Z(\s13.SbusIn [22]) );
  CNR2X1 U8751 ( .A(n4258), .B(n4194), .Z(\s13.SbusIn [49]) );
  CNR2X1 U8752 ( .A(n4259), .B(n4244), .Z(\s13.addr [59]) );
  CIVX2 U8753 ( .A(n4180), .Z(n4245) );
  CNR2X1 U8754 ( .A(n4259), .B(n4245), .Z(\s13.SbusIn [18]) );
  CNR2X1 U8755 ( .A(n4317), .B(n4236), .Z(\s0.addr [30]) );
  CNR2X1 U8756 ( .A(n4327), .B(n4246), .Z(\s0.addr [27]) );
  CIVDX4 U8757 ( .A(n4188), .Z0(n4314), .Z1(\s0.addr [12]) );
  CNR2X1 U8758 ( .A(n4314), .B(n4248), .Z(\s0.SbusIn [26]) );
  CNR2X1 U8759 ( .A(n4327), .B(n4230), .Z(\s0.addr [22]) );
  CIVDX4 U8760 ( .A(n4188), .Z0(n4321), .Z1(n3975) );
  CNR2X1 U8761 ( .A(n4321), .B(n4181), .Z(\s0.SbusIn [25]) );
  CNR2X1 U8762 ( .A(n4314), .B(n4182), .Z(\s0.addr [29]) );
  CIVDX4 U8763 ( .A(n4188), .Z0(n4307), .Z1(\s0.addr [13]) );
  CNR2X1 U8764 ( .A(n4307), .B(n4194), .Z(\s0.SbusIn [49]) );
  CNR2X1 U8765 ( .A(n4321), .B(n4249), .Z(\s0.SbusIn [50]) );
  CIVDX4 U8766 ( .A(n4188), .Z0(n4309), .Z1(n3940) );
  CNR2X1 U8767 ( .A(n4309), .B(n4183), .Z(\s0.SbusIn [10]) );
  CNR2X1 U8768 ( .A(n4319), .B(n4231), .Z(\s0.SbusIn [22]) );
  CIVDX4 U8769 ( .A(n4188), .Z0(n4311), .Z1(\s0.en ) );
  CNR2X1 U8770 ( .A(n4311), .B(n4184), .Z(\s0.addr [21]) );
  CNR2X1 U8771 ( .A(n4319), .B(n4252), .Z(\s0.addr [54]) );
  CIVX2 U8772 ( .A(n4185), .Z(n4198) );
  CNR2X1 U8773 ( .A(n4325), .B(n4198), .Z(\s0.SbusIn [0]) );
  CNR2X1 U8774 ( .A(n4309), .B(n4235), .Z(\s0.SbusIn [60]) );
  CNR2X1 U8775 ( .A(n4307), .B(n4186), .Z(\s0.addr [47]) );
  CNR2X1 U8776 ( .A(n4309), .B(n4187), .Z(\s0.SbusIn [6]) );
  CNR2X1 U8777 ( .A(n4319), .B(n4239), .Z(\s0.addr [53]) );
  CIVDX4 U8778 ( .A(n4188), .Z0(n4323), .Z1(n4106) );
  CNR2X1 U8779 ( .A(n4323), .B(n4189), .Z(\s0.addr [46]) );
  CIVX2 U8780 ( .A(n4190), .Z(n4241) );
  CNR2X1 U8781 ( .A(n4311), .B(n4241), .Z(\s0.SbusIn [1]) );
  CNR2X1 U8782 ( .A(n4325), .B(n4191), .Z(\s0.SbusIn [61]) );
  CIVX2 U8783 ( .A(n4192), .Z(n4214) );
  CNR2X1 U8784 ( .A(n4258), .B(n4214), .Z(\s13.SbusIn [2]) );
  CNR2X1 U8785 ( .A(n4259), .B(n4222), .Z(\s13.SbusIn [19]) );
  CNR2X1 U8786 ( .A(n4259), .B(n4241), .Z(\s13.SbusIn [1]) );
  CNR2X1 U8787 ( .A(n4259), .B(n4198), .Z(\s13.SbusIn [0]) );
  CIVX2 U8788 ( .A(n4193), .Z(n4282) );
  CNR2X1 U8789 ( .A(n4258), .B(n4282), .Z(\s13.SbusIn [9]) );
  CNR2X1 U8790 ( .A(n4258), .B(n4219), .Z(\s13.SbusIn [59]) );
  CNR2X1 U8791 ( .A(n4259), .B(n4206), .Z(\s13.addr [23]) );
  CNR2X1 U8792 ( .A(n4256), .B(n4194), .Z(\s2.SbusIn [49]) );
  CIVX2 U8793 ( .A(n4328), .Z(n4270) );
  CNR2X1 U8794 ( .A(n4255), .B(n4270), .Z(\s2.addr [25]) );
  CIVX2 U8795 ( .A(n4195), .Z(n4224) );
  CNR2X1 U8796 ( .A(n4255), .B(n4224), .Z(\s2.addr [26]) );
  CNR2X1 U8797 ( .A(n4256), .B(n4271), .Z(\s2.SbusIn [53]) );
  CIVX1 U8798 ( .A(n4196), .Z(n4315) );
  CNR2X1 U8799 ( .A(n4256), .B(n4315), .Z(\s2.SbusIn [37]) );
  CNR2X1 U8800 ( .A(n4256), .B(n4294), .Z(\s2.SbusIn [57]) );
  CNR2X1 U8801 ( .A(n4256), .B(n4227), .Z(\s2.SbusIn [21]) );
  CIVX2 U8802 ( .A(n4197), .Z(n4266) );
  CNR2X1 U8803 ( .A(n4255), .B(n4266), .Z(\s2.SbusIn [29]) );
  CNR2X1 U8804 ( .A(n4255), .B(n4310), .Z(\s2.SbusIn [17]) );
  CNR2X1 U8805 ( .A(n4256), .B(n4324), .Z(\s2.addr [44]) );
  CNR2X1 U8806 ( .A(n4256), .B(n4287), .Z(\s2.addr [32]) );
  CNR2X1 U8807 ( .A(n4255), .B(n4298), .Z(\s2.SbusIn [32]) );
  CNR2X1 U8808 ( .A(n4256), .B(n4272), .Z(\s2.addr [0]) );
  CNR2X1 U8809 ( .A(n4256), .B(n4198), .Z(\s2.SbusIn [0]) );
  CIVX2 U8810 ( .A(n4199), .Z(n4278) );
  CNR2X1 U8811 ( .A(n4255), .B(n4278), .Z(\s2.addr [24]) );
  CNR2X1 U8812 ( .A(n4256), .B(n4282), .Z(\s2.SbusIn [9]) );
  CIVX2 U8813 ( .A(n4200), .Z(n4277) );
  CNR2X1 U8814 ( .A(n4255), .B(n4277), .Z(\s2.SbusIn [3]) );
  CIVX2 U8815 ( .A(n4201), .Z(n4208) );
  CNR2X1 U8816 ( .A(n4255), .B(n4208), .Z(\s2.addr [55]) );
  CNR2X1 U8817 ( .A(n4255), .B(n4225), .Z(\s2.SbusIn [14]) );
  CNR2X1 U8818 ( .A(n4255), .B(n4285), .Z(\s2.addr [37]) );
  CNR2X1 U8819 ( .A(n4256), .B(n4276), .Z(\s2.addr [52]) );
  CIVX2 U8820 ( .A(n4202), .Z(n4301) );
  CNR2X1 U8821 ( .A(n4256), .B(n4301), .Z(\s2.addr [58]) );
  CNR2X1 U8822 ( .A(n4259), .B(n4300), .Z(\s13.addr [41]) );
  CNR2X1 U8823 ( .A(n4319), .B(n4214), .Z(\s0.SbusIn [2]) );
  CNR2X1 U8824 ( .A(n4258), .B(n4268), .Z(\s13.SbusIn [7]) );
  CNR2X1 U8825 ( .A(n4323), .B(n4203), .Z(\s0.addr [48]) );
  CIVX2 U8826 ( .A(n4204), .Z(n4281) );
  CNR2X1 U8827 ( .A(n4258), .B(n4281), .Z(\s13.addr [38]) );
  CNR2X1 U8828 ( .A(n4317), .B(n4208), .Z(\s0.addr [55]) );
  CNR2X1 U8829 ( .A(n4314), .B(n4205), .Z(\s0.addr [20]) );
  CNR2X1 U8830 ( .A(n4259), .B(n4292), .Z(\s13.SbusIn [31]) );
  CNR2X1 U8831 ( .A(n4309), .B(n4206), .Z(\s0.addr [23]) );
  CNR2X1 U8832 ( .A(n4259), .B(n4210), .Z(\s13.SbusIn [23]) );
  CIVX2 U8833 ( .A(n4207), .Z(n4291) );
  CNR2X1 U8834 ( .A(n4258), .B(n4291), .Z(\s13.addr [57]) );
  CNR2X1 U8835 ( .A(n4258), .B(n4208), .Z(\s13.addr [55]) );
  CNR2X1 U8836 ( .A(n4319), .B(n4209), .Z(\s0.SbusIn [11]) );
  CNR2X1 U8837 ( .A(n4323), .B(n4233), .Z(\s0.SbusIn [51]) );
  CNR2X1 U8838 ( .A(n4317), .B(n4210), .Z(\s0.SbusIn [23]) );
  CNR2X1 U8839 ( .A(n4259), .B(n4224), .Z(\s13.addr [26]) );
  CNR2X1 U8840 ( .A(n4321), .B(n4211), .Z(\s0.SbusIn [62]) );
  CNR2X1 U8841 ( .A(n4307), .B(n4213), .Z(\s0.SbusIn [52]) );
  CNR2X1 U8842 ( .A(n4259), .B(n4302), .Z(\s13.SbusIn [12]) );
  CNR2X1 U8843 ( .A(n4311), .B(n4212), .Z(\s0.SbusIn [27]) );
  CNR2X1 U8844 ( .A(n4258), .B(n4301), .Z(\s13.addr [58]) );
  CNR2X1 U8845 ( .A(n4258), .B(n4270), .Z(\s13.addr [25]) );
  CNR2X1 U8846 ( .A(n4259), .B(n4296), .Z(\s13.addr [61]) );
  CNR2X1 U8847 ( .A(n4256), .B(n4288), .Z(\s2.SbusIn [16]) );
  CNR2X1 U8848 ( .A(n4255), .B(n4291), .Z(\s2.addr [57]) );
  CNR2X1 U8849 ( .A(n4255), .B(n4283), .Z(\s2.SbusIn [56]) );
  CNR2X1 U8850 ( .A(n4255), .B(n4213), .Z(\s2.SbusIn [52]) );
  CNR2X1 U8851 ( .A(n4256), .B(n4214), .Z(\s2.SbusIn [2]) );
  CNR2X1 U8852 ( .A(n4256), .B(n4305), .Z(\s2.addr [31]) );
  CNR2X1 U8853 ( .A(n4255), .B(n4264), .Z(\s2.addr [51]) );
  CNR2X1 U8854 ( .A(n4256), .B(n4220), .Z(\s2.SbusIn [34]) );
  CNR2X1 U8855 ( .A(n4255), .B(n4267), .Z(\s2.addr [39]) );
  CNR2X1 U8856 ( .A(n4255), .B(n4216), .Z(\s2.addr [35]) );
  CIVDX1 U8857 ( .A(n4215), .Z0(n4279), .Z1(n3376) );
  CNR2X1 U8858 ( .A(n4256), .B(n4279), .Z(\s2.SbusIn [36]) );
  CNR2X1 U8859 ( .A(n4323), .B(n4216), .Z(\s0.addr [35]) );
  CNR2X1 U8860 ( .A(n4317), .B(n4217), .Z(\s0.addr [28]) );
  CNR2X1 U8861 ( .A(n4323), .B(n4218), .Z(\s0.SbusIn [47]) );
  CNR2X1 U8862 ( .A(n4309), .B(n4219), .Z(\s0.SbusIn [59]) );
  CNR2X1 U8863 ( .A(n4325), .B(n4220), .Z(\s0.SbusIn [34]) );
  CNR2X1 U8864 ( .A(n4327), .B(n4240), .Z(\s0.SbusIn [33]) );
  CNR2X1 U8865 ( .A(n4321), .B(n4221), .Z(\s0.addr [34]) );
  CNR2X1 U8866 ( .A(n4327), .B(n4222), .Z(\s0.SbusIn [19]) );
  CNR2X1 U8867 ( .A(n4321), .B(n4251), .Z(\s0.addr [60]) );
  CNR2X1 U8868 ( .A(n4309), .B(n4223), .Z(\s0.addr [42]) );
  CNR2X1 U8869 ( .A(n4309), .B(n4224), .Z(\s0.addr [26]) );
  CNR2X1 U8870 ( .A(n4319), .B(n4244), .Z(\s0.addr [59]) );
  CNR2X1 U8871 ( .A(n4319), .B(n4225), .Z(\s0.SbusIn [14]) );
  CNR2X1 U8872 ( .A(n4323), .B(n4247), .Z(\s0.SbusIn [13]) );
  CNR2X1 U8873 ( .A(n4314), .B(n4226), .Z(\s0.SbusIn [48]) );
  CNR2X1 U8874 ( .A(n4314), .B(n4245), .Z(\s0.SbusIn [18]) );
  CNR2X1 U8875 ( .A(n4307), .B(n4227), .Z(\s0.SbusIn [21]) );
  CNR2X1 U8876 ( .A(n4307), .B(n4228), .Z(\s0.SbusIn [5]) );
  CNR2X1 U8877 ( .A(n4311), .B(n4238), .Z(\s0.addr [45]) );
  CNR2X1 U8878 ( .A(n4311), .B(n4229), .Z(\s0.addr [63]) );
  CNR2X1 U8879 ( .A(n4325), .B(n4234), .Z(\s0.SbusIn [58]) );
  CNR2X1 U8880 ( .A(n4259), .B(n4230), .Z(\s13.addr [22]) );
  CNR2X1 U8881 ( .A(n4259), .B(n4266), .Z(\s13.SbusIn [29]) );
  CNR2X1 U8882 ( .A(n4256), .B(n4231), .Z(\s2.SbusIn [22]) );
  CIVDX1 U8883 ( .A(n4232), .Z0(n4290), .Z1(n3331) );
  CNR2X1 U8884 ( .A(n4255), .B(n4290), .Z(\s2.SbusIn [38]) );
  CNR2X1 U8885 ( .A(n4255), .B(n4233), .Z(\s2.SbusIn [51]) );
  CNR2X1 U8886 ( .A(n4256), .B(n4263), .Z(\s2.SbusIn [54]) );
  CNR2X1 U8887 ( .A(n4256), .B(n4308), .Z(\s2.SbusIn [55]) );
  CNR2X1 U8888 ( .A(n4256), .B(n4234), .Z(\s2.SbusIn [58]) );
  CNR2X1 U8889 ( .A(n4255), .B(n4235), .Z(\s2.SbusIn [60]) );
  CNR2X1 U8890 ( .A(n4256), .B(n4318), .Z(\s2.addr [2]) );
  CNR2X1 U8891 ( .A(n4255), .B(n4246), .Z(\s2.addr [27]) );
  CNR2X1 U8892 ( .A(n4256), .B(n4236), .Z(\s2.addr [30]) );
  CIVX2 U8893 ( .A(n4237), .Z(n4274) );
  CNR2X1 U8894 ( .A(n4256), .B(n4274), .Z(\s2.SbusIn [35]) );
  CNR2X1 U8895 ( .A(n4255), .B(n4306), .Z(\s2.addr [33]) );
  CNR2X1 U8896 ( .A(n4255), .B(n4281), .Z(\s2.addr [38]) );
  CNR2X1 U8897 ( .A(n4255), .B(n4238), .Z(\s2.addr [45]) );
  CNR2X1 U8898 ( .A(n4255), .B(n4260), .Z(\s2.addr [50]) );
  CNR2X1 U8899 ( .A(n4255), .B(n4239), .Z(\s2.addr [53]) );
  CNR2X1 U8900 ( .A(n4256), .B(n4240), .Z(\s2.SbusIn [33]) );
  CNR2X1 U8901 ( .A(n4256), .B(n4241), .Z(\s2.SbusIn [1]) );
  CIVX2 U8902 ( .A(n4242), .Z(n4313) );
  CNR2X1 U8903 ( .A(n4255), .B(n4313), .Z(\s2.addr [56]) );
  CIVX2 U8904 ( .A(n4243), .Z(n4262) );
  CNR2X1 U8905 ( .A(n4256), .B(n4262), .Z(\s2.SbusIn [4]) );
  CNR2X1 U8906 ( .A(n4256), .B(n4244), .Z(\s2.addr [59]) );
  CNR2X1 U8907 ( .A(n4256), .B(n4251), .Z(\s2.addr [60]) );
  CNR2X1 U8908 ( .A(n4256), .B(n4297), .Z(\s2.SbusIn [15]) );
  CNR2X1 U8909 ( .A(n4255), .B(n4245), .Z(\s2.SbusIn [18]) );
  CNR2X1 U8910 ( .A(n4258), .B(n4246), .Z(\s13.addr [27]) );
  CNR2X1 U8911 ( .A(n4258), .B(n4316), .Z(\s13.SbusIn [8]) );
  CNR2X1 U8912 ( .A(n4259), .B(n4247), .Z(\s13.SbusIn [13]) );
  CNR2X1 U8913 ( .A(n4259), .B(n4278), .Z(\s13.addr [24]) );
  CNR2X1 U8914 ( .A(n4258), .B(n4248), .Z(\s13.SbusIn [26]) );
  CNR2X1 U8915 ( .A(n4258), .B(n4249), .Z(\s13.SbusIn [50]) );
  CNR2X1 U8916 ( .A(n4259), .B(n4313), .Z(\s13.addr [56]) );
  CNR2X1 U8917 ( .A(n4259), .B(n4250), .Z(\s13.addr [62]) );
  CNR2X1 U8918 ( .A(n4258), .B(n4275), .Z(\s13.addr [49]) );
  CNR2X1 U8919 ( .A(n4258), .B(n4251), .Z(\s13.addr [60]) );
  CNR2X1 U8920 ( .A(n4259), .B(n4295), .Z(\s13.SbusIn [20]) );
  CNR2X1 U8921 ( .A(n4259), .B(n4252), .Z(\s13.addr [54]) );
  CNR2X1 U8922 ( .A(n4258), .B(n4280), .Z(\s13.SbusIn [24]) );
  CNR2X1 U8923 ( .A(n4259), .B(n4262), .Z(\s13.SbusIn [4]) );
  CNR2X1 U8924 ( .A(n4258), .B(n4277), .Z(\s13.SbusIn [3]) );
  CNR2X1 U8925 ( .A(n4255), .B(n4253), .Z(\s2.addr [5]) );
  CNR2X1 U8926 ( .A(n4255), .B(n4254), .Z(\s2.addr [4]) );
  CNR2X1 U8927 ( .A(n4256), .B(n4326), .Z(\s2.addr [6]) );
  CNR2X1 U8928 ( .A(n4258), .B(n4257), .Z(\s13.addr [7]) );
  CNR2X1 U8929 ( .A(n4259), .B(n4293), .Z(\s13.SbusIn [39]) );
  CNR2X1 U8930 ( .A(n4321), .B(n4260), .Z(\s0.addr [50]) );
  CNR2X1 U8931 ( .A(n4311), .B(n4261), .Z(\s0.SbusIn [63]) );
  CNR2X1 U8932 ( .A(n4323), .B(n4262), .Z(\s0.SbusIn [4]) );
  CNR2X1 U8933 ( .A(n4317), .B(n4263), .Z(\s0.SbusIn [54]) );
  CNR2X1 U8934 ( .A(n4321), .B(n4264), .Z(\s0.addr [51]) );
  CNR2X1 U8935 ( .A(n4325), .B(n4265), .Z(\s0.SbusIn [40]) );
  CNR2X1 U8936 ( .A(n4317), .B(n4266), .Z(\s0.SbusIn [29]) );
  CNR2X1 U8937 ( .A(n4314), .B(n4267), .Z(\s0.addr [39]) );
  CNR2X1 U8938 ( .A(n4307), .B(n4268), .Z(\s0.SbusIn [7]) );
  CNR2X1 U8939 ( .A(n4323), .B(n4269), .Z(\s0.SbusIn [41]) );
  CNR2X1 U8940 ( .A(n4309), .B(n4270), .Z(\s0.addr [25]) );
  CNR2X1 U8941 ( .A(n4327), .B(n4271), .Z(\s0.SbusIn [53]) );
  CNR2X1 U8942 ( .A(n4314), .B(n4272), .Z(\s0.addr [0]) );
  CNR2X1 U8943 ( .A(n4321), .B(n4273), .Z(\s0.SbusIn [28]) );
  CNR2X1 U8944 ( .A(n4317), .B(n4274), .Z(\s0.SbusIn [35]) );
  CNR2X1 U8945 ( .A(n4309), .B(n4275), .Z(\s0.addr [49]) );
  CNR2X1 U8946 ( .A(n4319), .B(n4276), .Z(\s0.addr [52]) );
  CNR2X1 U8947 ( .A(n4307), .B(n4277), .Z(\s0.SbusIn [3]) );
  CNR2X1 U8948 ( .A(n4311), .B(n4278), .Z(\s0.addr [24]) );
  CNR2X1 U8949 ( .A(n4323), .B(n4279), .Z(\s0.SbusIn [36]) );
  CNR2X1 U8950 ( .A(n4325), .B(n4280), .Z(\s0.SbusIn [24]) );
  CNR2X1 U8951 ( .A(n4327), .B(n4281), .Z(\s0.addr [38]) );
  CNR2X1 U8952 ( .A(n4317), .B(n4282), .Z(\s0.SbusIn [9]) );
  CNR2X1 U8953 ( .A(n4314), .B(n4283), .Z(\s0.SbusIn [56]) );
  CNR2X1 U8954 ( .A(n4307), .B(n4284), .Z(\s0.addr [43]) );
  CNR2X1 U8955 ( .A(n4311), .B(n4285), .Z(\s0.addr [37]) );
  CNR2X1 U8956 ( .A(n4325), .B(n4286), .Z(\s0.SbusIn [43]) );
  CNR2X1 U8957 ( .A(n4321), .B(n4287), .Z(\s0.addr [32]) );
  CNR2X1 U8958 ( .A(n4314), .B(n4288), .Z(\s0.SbusIn [16]) );
  CNR2X1 U8959 ( .A(n4307), .B(n4289), .Z(\s0.SbusIn [46]) );
  CNR2X1 U8960 ( .A(n4311), .B(n4290), .Z(\s0.SbusIn [38]) );
  CNR2X1 U8961 ( .A(n4327), .B(n4291), .Z(\s0.addr [57]) );
  CNR2X1 U8962 ( .A(n4325), .B(n4292), .Z(\s0.SbusIn [31]) );
  CNR2X1 U8963 ( .A(n4319), .B(n4293), .Z(\s0.SbusIn [39]) );
  CNR2X1 U8964 ( .A(n4314), .B(n4294), .Z(\s0.SbusIn [57]) );
  CNR2X1 U8965 ( .A(n4307), .B(n4295), .Z(\s0.SbusIn [20]) );
  CNR2X1 U8966 ( .A(n4327), .B(n4296), .Z(\s0.addr [61]) );
  CNR2X1 U8967 ( .A(n4321), .B(n4297), .Z(\s0.SbusIn [15]) );
  CNR2X1 U8968 ( .A(n4311), .B(n4298), .Z(\s0.SbusIn [32]) );
  CNR2X1 U8969 ( .A(n4309), .B(n4299), .Z(\s0.SbusIn [42]) );
  CNR2X1 U8970 ( .A(n4323), .B(n4300), .Z(\s0.addr [41]) );
  CNR2X1 U8971 ( .A(n4325), .B(n4301), .Z(\s0.addr [58]) );
  CNR2X1 U8972 ( .A(n4327), .B(n4302), .Z(\s0.SbusIn [12]) );
  CNR2X1 U8973 ( .A(n4317), .B(n4303), .Z(\s0.SbusIn [45]) );
  CNR2X1 U8974 ( .A(n4309), .B(n4304), .Z(\s0.SbusIn [30]) );
  CNR2X1 U8975 ( .A(n4321), .B(n4305), .Z(\s0.addr [31]) );
  CNR2X1 U8976 ( .A(n4307), .B(n4306), .Z(\s0.addr [33]) );
  CNR2X1 U8977 ( .A(n4309), .B(n4308), .Z(\s0.SbusIn [55]) );
  CNR2X1 U8978 ( .A(n4311), .B(n4310), .Z(\s0.SbusIn [17]) );
  CNR2X1 U8979 ( .A(n4319), .B(n4312), .Z(\s0.addr [40]) );
  CNR2X1 U8980 ( .A(n4314), .B(n4313), .Z(\s0.addr [56]) );
  CNR2X1 U8981 ( .A(n4323), .B(n4315), .Z(\s0.SbusIn [37]) );
  CNR2X1 U8982 ( .A(n4317), .B(n4316), .Z(\s0.SbusIn [8]) );
  CNR2X1 U8983 ( .A(n4319), .B(n4318), .Z(\s0.addr [2]) );
  CNR2X1 U8984 ( .A(n4321), .B(n4320), .Z(\s0.SbusIn [44]) );
  CNR2X1 U8985 ( .A(n4323), .B(n4322), .Z(\s0.addr [36]) );
  CNR2X1 U8986 ( .A(n4325), .B(n4324), .Z(\s0.addr [44]) );
  CNR2X1 U8987 ( .A(n4327), .B(n4326), .Z(\s0.addr [6]) );
  CAN2X1 U8988 ( .A(\s9.en ), .B(n4328), .Z(\s9.addr [25]) );
  CAN2X1 U8989 ( .A(\s12.addr[11] ), .B(n3456), .Z(\s12.addr [7]) );
  CAN2XL U8990 ( .A(n4405), .B(n4333), .Z(\s5.addr [3]) );
  CAN2XL U8991 ( .A(\s6.en ), .B(n4333), .Z(\s6.addr [3]) );
  CAN2XL U8992 ( .A(\s14.addr[18] ), .B(n4333), .Z(\s14.addr [3]) );
  CAN2XL U8993 ( .A(\s4.addr [19]), .B(n4337), .Z(\s4.addr [0]) );
  CAN2XL U8994 ( .A(n4405), .B(n4337), .Z(\s5.addr [0]) );
  CAN2XL U8995 ( .A(n1844), .B(n4339), .Z(\s5.addr [1]) );
  CAN2XL U8996 ( .A(\s3.addr [18]), .B(n4337), .Z(\s3.addr [0]) );
  CAN2XL U8997 ( .A(\s3.addr[14] ), .B(n4339), .Z(\s3.addr [1]) );
  CAN2XL U8998 ( .A(\s14.addr[17] ), .B(n4337), .Z(\s14.addr [0]) );
  CAN2XL U8999 ( .A(\s14.addr [11]), .B(n4338), .Z(\s14.addr [4]) );
  CAN2XL U9000 ( .A(\s12.addr[11] ), .B(n4337), .Z(\s12.addr [0]) );
  CAN2XL U9001 ( .A(\s12.addr[16] ), .B(n4330), .Z(\s12.addr [2]) );
  CAN2XL U9002 ( .A(\s12.addr[16] ), .B(n4334), .Z(\s12.addr [4]) );
  CAN2XL U9003 ( .A(\s12.addr[10] ), .B(n4331), .Z(\s12.addr [20]) );
  CAN2XL U9004 ( .A(n4332), .B(n4337), .Z(\s11.addr [0]) );
  CAN2XL U9005 ( .A(\s10.en ), .B(n4337), .Z(\s10.addr [0]) );
  CAN2XL U9006 ( .A(\s10.en ), .B(n4339), .Z(\s10.addr [1]) );
  CAN2XL U9007 ( .A(\s10.en ), .B(n4333), .Z(\s10.addr [3]) );
  CAN2XL U9008 ( .A(\s10.en ), .B(n4334), .Z(\s10.addr [4]) );
  CAN2XL U9009 ( .A(\s10.en ), .B(n4335), .Z(\s10.addr [8]) );
  CAN2XL U9010 ( .A(\s9.addr[7] ), .B(n4337), .Z(\s9.addr [0]) );
  CAN2XL U9011 ( .A(\s8.addr[17] ), .B(n4337), .Z(\s8.addr [0]) );
  CAN2XL U9012 ( .A(\s8.addr[15] ), .B(n4339), .Z(\s8.addr [1]) );
  CAN2XL U9013 ( .A(\s8.addr[17] ), .B(n4338), .Z(\s8.addr [4]) );
  CAN2XL U9014 ( .A(\s8.addr[17] ), .B(n4335), .Z(\s8.addr [8]) );
  CAN2XL U9015 ( .A(n4336), .B(n4337), .Z(\s7.addr [0]) );
  CAN2XL U9016 ( .A(n4336), .B(n4338), .Z(\s7.addr [4]) );
  CAN2XL U9017 ( .A(\s6.addr [17]), .B(n4337), .Z(\s6.addr [0]) );
  CAN2XL U9018 ( .A(\s6.addr [17]), .B(n4339), .Z(\s6.addr [1]) );
  CAN2XL U9019 ( .A(\s6.en ), .B(n4338), .Z(\s6.addr [4]) );
  CAN2XL U9020 ( .A(n5445), .B(n4338), .Z(\s5.addr [4]) );
  CAN2XL U9021 ( .A(\s4.en ), .B(n4339), .Z(\s4.addr [1]) );
endmodule

